VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mac_cluster
  CLASS BLOCK ;
  FOREIGN mac_cluster ;
  ORIGIN 0.000 0.000 ;
  SIZE 497.345 BY 508.065 ;
  PIN A0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.930 504.065 186.210 508.065 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 272.040 497.345 272.640 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 418.690 504.065 418.970 508.065 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.650 504.065 200.930 508.065 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END A0[7]
  PIN A1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 175.810 504.065 176.090 508.065 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 466.520 497.345 467.120 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 261.370 504.065 261.650 508.065 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 287.130 504.065 287.410 508.065 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 504.065 18.770 508.065 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.490 504.065 271.770 508.065 ;
    END
  END A1[7]
  PIN A2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 449.050 504.065 449.330 508.065 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END A2[6]
  PIN A2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 443.400 497.345 444.000 ;
    END
  END A2[7]
  PIN A3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.530 504.065 236.810 508.065 ;
    END
  END A3[0]
  PIN A3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END A3[1]
  PIN A3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 463.770 504.065 464.050 508.065 ;
    END
  END A3[2]
  PIN A3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.170 504.065 206.450 508.065 ;
    END
  END A3[3]
  PIN A3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END A3[4]
  PIN A3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END A3[5]
  PIN A3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END A3[6]
  PIN A3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.090 504.065 69.370 508.065 ;
    END
  END A3[7]
  PIN B0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END B0[0]
  PIN B0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END B0[1]
  PIN B0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END B0[2]
  PIN B0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END B0[3]
  PIN B0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 219.000 497.345 219.600 ;
    END
  END B0[4]
  PIN B0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 226.410 504.065 226.690 508.065 ;
    END
  END B0[5]
  PIN B0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 504.065 73.970 508.065 ;
    END
  END B0[6]
  PIN B0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END B0[7]
  PIN B1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.450 504.065 145.730 508.065 ;
    END
  END B1[0]
  PIN B1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 368.600 497.345 369.200 ;
    END
  END B1[1]
  PIN B1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 152.360 497.345 152.960 ;
    END
  END B1[2]
  PIN B1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END B1[3]
  PIN B1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.690 504.065 372.970 508.065 ;
    END
  END B1[4]
  PIN B1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END B1[5]
  PIN B1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.570 504.065 155.850 508.065 ;
    END
  END B1[6]
  PIN B1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 242.120 497.345 242.720 ;
    END
  END B1[7]
  PIN B2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END B2[0]
  PIN B2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END B2[1]
  PIN B2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END B2[2]
  PIN B2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 114.280 497.345 114.880 ;
    END
  END B2[3]
  PIN B2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.170 504.065 160.450 508.065 ;
    END
  END B2[4]
  PIN B2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 504.065 23.370 508.065 ;
    END
  END B2[5]
  PIN B2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END B2[6]
  PIN B2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 278.840 497.345 279.440 ;
    END
  END B2[7]
  PIN B3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 77.560 497.345 78.160 ;
    END
  END B3[0]
  PIN B3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END B3[1]
  PIN B3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END B3[2]
  PIN B3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 481.480 497.345 482.080 ;
    END
  END B3[3]
  PIN B3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 212.200 497.345 212.800 ;
    END
  END B3[4]
  PIN B3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 504.065 28.890 508.065 ;
    END
  END B3[5]
  PIN B3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END B3[6]
  PIN B3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 107.480 497.345 108.080 ;
    END
  END B3[7]
  PIN cfg[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.770 504.065 257.050 508.065 ;
    END
  END cfg[0]
  PIN cfg[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END cfg[100]
  PIN cfg[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END cfg[101]
  PIN cfg[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END cfg[102]
  PIN cfg[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 504.065 49.130 508.065 ;
    END
  END cfg[103]
  PIN cfg[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END cfg[104]
  PIN cfg[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END cfg[105]
  PIN cfg[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 428.440 497.345 429.040 ;
    END
  END cfg[106]
  PIN cfg[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END cfg[107]
  PIN cfg[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END cfg[108]
  PIN cfg[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.570 504.065 109.850 508.065 ;
    END
  END cfg[109]
  PIN cfg[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END cfg[10]
  PIN cfg[110]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END cfg[110]
  PIN cfg[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END cfg[111]
  PIN cfg[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END cfg[112]
  PIN cfg[113]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 204.040 497.345 204.640 ;
    END
  END cfg[113]
  PIN cfg[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 248.920 497.345 249.520 ;
    END
  END cfg[114]
  PIN cfg[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.330 504.065 89.610 508.065 ;
    END
  END cfg[115]
  PIN cfg[116]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END cfg[116]
  PIN cfg[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 428.810 504.065 429.090 508.065 ;
    END
  END cfg[117]
  PIN cfg[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END cfg[118]
  PIN cfg[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END cfg[119]
  PIN cfg[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END cfg[11]
  PIN cfg[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.690 504.065 119.970 508.065 ;
    END
  END cfg[120]
  PIN cfg[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 24.520 497.345 25.120 ;
    END
  END cfg[121]
  PIN cfg[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END cfg[122]
  PIN cfg[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END cfg[123]
  PIN cfg[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 361.800 497.345 362.400 ;
    END
  END cfg[124]
  PIN cfg[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 504.065 33.490 508.065 ;
    END
  END cfg[125]
  PIN cfg[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 257.080 497.345 257.680 ;
    END
  END cfg[126]
  PIN cfg[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END cfg[127]
  PIN cfg[128]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END cfg[128]
  PIN cfg[129]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END cfg[129]
  PIN cfg[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END cfg[12]
  PIN cfg[130]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END cfg[130]
  PIN cfg[131]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.850 504.065 348.130 508.065 ;
    END
  END cfg[131]
  PIN cfg[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.090 504.065 322.370 508.065 ;
    END
  END cfg[13]
  PIN cfg[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END cfg[14]
  PIN cfg[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END cfg[15]
  PIN cfg[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END cfg[16]
  PIN cfg[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 291.730 504.065 292.010 508.065 ;
    END
  END cfg[17]
  PIN cfg[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 353.640 497.345 354.240 ;
    END
  END cfg[18]
  PIN cfg[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END cfg[19]
  PIN cfg[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END cfg[1]
  PIN cfg[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.770 504.065 211.050 508.065 ;
    END
  END cfg[20]
  PIN cfg[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 92.520 497.345 93.120 ;
    END
  END cfg[21]
  PIN cfg[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 174.120 497.345 174.720 ;
    END
  END cfg[22]
  PIN cfg[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END cfg[23]
  PIN cfg[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 17.720 497.345 18.320 ;
    END
  END cfg[24]
  PIN cfg[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END cfg[25]
  PIN cfg[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END cfg[26]
  PIN cfg[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.730 504.065 338.010 508.065 ;
    END
  END cfg[27]
  PIN cfg[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 433.410 504.065 433.690 508.065 ;
    END
  END cfg[28]
  PIN cfg[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END cfg[29]
  PIN cfg[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END cfg[2]
  PIN cfg[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END cfg[30]
  PIN cfg[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 316.920 497.345 317.520 ;
    END
  END cfg[31]
  PIN cfg[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 469.290 504.065 469.570 508.065 ;
    END
  END cfg[32]
  PIN cfg[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 251.250 504.065 251.530 508.065 ;
    END
  END cfg[33]
  PIN cfg[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END cfg[34]
  PIN cfg[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END cfg[35]
  PIN cfg[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END cfg[36]
  PIN cfg[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END cfg[37]
  PIN cfg[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 54.440 497.345 55.040 ;
    END
  END cfg[38]
  PIN cfg[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 383.560 497.345 384.160 ;
    END
  END cfg[39]
  PIN cfg[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 458.360 497.345 458.960 ;
    END
  END cfg[3]
  PIN cfg[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END cfg[40]
  PIN cfg[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.730 504.065 85.010 508.065 ;
    END
  END cfg[41]
  PIN cfg[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END cfg[42]
  PIN cfg[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END cfg[43]
  PIN cfg[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 129.240 497.345 129.840 ;
    END
  END cfg[44]
  PIN cfg[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END cfg[45]
  PIN cfg[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 406.680 497.345 407.280 ;
    END
  END cfg[46]
  PIN cfg[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 398.450 504.065 398.730 508.065 ;
    END
  END cfg[47]
  PIN cfg[48]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END cfg[48]
  PIN cfg[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 504.065 79.490 508.065 ;
    END
  END cfg[49]
  PIN cfg[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 504.065 170.570 508.065 ;
    END
  END cfg[4]
  PIN cfg[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END cfg[50]
  PIN cfg[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 459.170 504.065 459.450 508.065 ;
    END
  END cfg[51]
  PIN cfg[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END cfg[52]
  PIN cfg[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END cfg[53]
  PIN cfg[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END cfg[54]
  PIN cfg[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END cfg[55]
  PIN cfg[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END cfg[56]
  PIN cfg[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END cfg[57]
  PIN cfg[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 382.810 504.065 383.090 508.065 ;
    END
  END cfg[58]
  PIN cfg[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END cfg[59]
  PIN cfg[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 388.330 504.065 388.610 508.065 ;
    END
  END cfg[5]
  PIN cfg[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 488.280 497.345 488.880 ;
    END
  END cfg[60]
  PIN cfg[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 293.800 497.345 294.400 ;
    END
  END cfg[61]
  PIN cfg[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 297.250 504.065 297.530 508.065 ;
    END
  END cfg[62]
  PIN cfg[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 144.200 497.345 144.800 ;
    END
  END cfg[63]
  PIN cfg[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END cfg[64]
  PIN cfg[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END cfg[65]
  PIN cfg[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 504.065 105.250 508.065 ;
    END
  END cfg[66]
  PIN cfg[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 504.065 3.130 508.065 ;
    END
  END cfg[67]
  PIN cfg[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END cfg[68]
  PIN cfg[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END cfg[69]
  PIN cfg[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 301.850 504.065 302.130 508.065 ;
    END
  END cfg[6]
  PIN cfg[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END cfg[70]
  PIN cfg[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 159.160 497.345 159.760 ;
    END
  END cfg[71]
  PIN cfg[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END cfg[72]
  PIN cfg[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END cfg[73]
  PIN cfg[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 165.690 504.065 165.970 508.065 ;
    END
  END cfg[74]
  PIN cfg[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END cfg[75]
  PIN cfg[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END cfg[76]
  PIN cfg[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END cfg[77]
  PIN cfg[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 32.680 497.345 33.280 ;
    END
  END cfg[78]
  PIN cfg[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.050 504.065 403.330 508.065 ;
    END
  END cfg[79]
  PIN cfg[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END cfg[7]
  PIN cfg[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END cfg[80]
  PIN cfg[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END cfg[81]
  PIN cfg[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END cfg[82]
  PIN cfg[83]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END cfg[83]
  PIN cfg[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 494.130 504.065 494.410 508.065 ;
    END
  END cfg[84]
  PIN cfg[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.970 504.065 358.250 508.065 ;
    END
  END cfg[85]
  PIN cfg[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.490 504.065 317.770 508.065 ;
    END
  END cfg[86]
  PIN cfg[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 197.240 497.345 197.840 ;
    END
  END cfg[87]
  PIN cfg[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 332.210 504.065 332.490 508.065 ;
    END
  END cfg[88]
  PIN cfg[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END cfg[89]
  PIN cfg[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 331.880 497.345 332.480 ;
    END
  END cfg[8]
  PIN cfg[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END cfg[90]
  PIN cfg[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END cfg[91]
  PIN cfg[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END cfg[92]
  PIN cfg[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END cfg[93]
  PIN cfg[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END cfg[94]
  PIN cfg[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 504.065 115.370 508.065 ;
    END
  END cfg[95]
  PIN cfg[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 99.320 497.345 99.920 ;
    END
  END cfg[96]
  PIN cfg[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END cfg[97]
  PIN cfg[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END cfg[98]
  PIN cfg[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END cfg[99]
  PIN cfg[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 413.480 497.345 414.080 ;
    END
  END cfg[9]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 473.890 504.065 474.170 508.065 ;
    END
  END clk
  PIN cset
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 493.345 227.160 497.345 227.760 ;
    END
  END cset
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 277.010 504.065 277.290 508.065 ;
    END
  END en
  PIN out0[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END out0[0]
  PIN out0[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.170 504.065 413.450 508.065 ;
    END
  END out0[10]
  PIN out0[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 263.880 497.345 264.480 ;
    END
  END out0[11]
  PIN out0[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 421.640 497.345 422.240 ;
    END
  END out0[12]
  PIN out0[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 301.960 497.345 302.560 ;
    END
  END out0[13]
  PIN out0[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 122.440 497.345 123.040 ;
    END
  END out0[14]
  PIN out0[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.410 504.065 180.690 508.065 ;
    END
  END out0[15]
  PIN out0[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.930 504.065 140.210 508.065 ;
    END
  END out0[16]
  PIN out0[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 125.210 504.065 125.490 508.065 ;
    END
  END out0[17]
  PIN out0[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END out0[18]
  PIN out0[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END out0[19]
  PIN out0[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 338.680 497.345 339.280 ;
    END
  END out0[1]
  PIN out0[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END out0[20]
  PIN out0[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END out0[21]
  PIN out0[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END out0[22]
  PIN out0[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END out0[23]
  PIN out0[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 220.890 504.065 221.170 508.065 ;
    END
  END out0[24]
  PIN out0[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 378.210 504.065 378.490 508.065 ;
    END
  END out0[25]
  PIN out0[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 398.520 497.345 399.120 ;
    END
  END out0[26]
  PIN out0[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 451.560 497.345 452.160 ;
    END
  END out0[27]
  PIN out0[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.450 504.065 53.730 508.065 ;
    END
  END out0[28]
  PIN out0[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 323.720 497.345 324.320 ;
    END
  END out0[29]
  PIN out0[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 453.650 504.065 453.930 508.065 ;
    END
  END out0[2]
  PIN out0[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END out0[30]
  PIN out0[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END out0[31]
  PIN out0[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END out0[3]
  PIN out0[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 39.480 497.345 40.080 ;
    END
  END out0[4]
  PIN out0[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 376.760 497.345 377.360 ;
    END
  END out0[5]
  PIN out0[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 342.330 504.065 342.610 508.065 ;
    END
  END out0[6]
  PIN out0[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 308.760 497.345 309.360 ;
    END
  END out0[7]
  PIN out0[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END out0[8]
  PIN out0[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.010 504.065 484.290 508.065 ;
    END
  END out0[9]
  PIN out1[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 327.610 504.065 327.890 508.065 ;
    END
  END out1[0]
  PIN out1[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 346.840 497.345 347.440 ;
    END
  END out1[10]
  PIN out1[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 436.600 497.345 437.200 ;
    END
  END out1[11]
  PIN out1[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END out1[12]
  PIN out1[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END out1[13]
  PIN out1[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.330 504.065 43.610 508.065 ;
    END
  END out1[14]
  PIN out1[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 307.370 504.065 307.650 508.065 ;
    END
  END out1[15]
  PIN out1[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END out1[16]
  PIN out1[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 189.080 497.345 189.680 ;
    END
  END out1[17]
  PIN out1[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.730 504.065 39.010 508.065 ;
    END
  END out1[18]
  PIN out1[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END out1[19]
  PIN out1[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END out1[1]
  PIN out1[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 473.320 497.345 473.920 ;
    END
  END out1[20]
  PIN out1[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.290 504.065 423.570 508.065 ;
    END
  END out1[21]
  PIN out1[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END out1[22]
  PIN out1[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END out1[23]
  PIN out1[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 504.065 130.090 508.065 ;
    END
  END out1[24]
  PIN out1[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END out1[25]
  PIN out1[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END out1[26]
  PIN out1[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 479.410 504.065 479.690 508.065 ;
    END
  END out1[27]
  PIN out1[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 167.320 497.345 167.920 ;
    END
  END out1[28]
  PIN out1[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.130 0.000 448.410 4.000 ;
    END
  END out1[29]
  PIN out1[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END out1[2]
  PIN out1[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END out1[30]
  PIN out1[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.970 504.065 13.250 508.065 ;
    END
  END out1[31]
  PIN out1[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 69.400 497.345 70.000 ;
    END
  END out1[3]
  PIN out1[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END out1[4]
  PIN out1[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END out1[5]
  PIN out1[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END out1[6]
  PIN out1[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 182.280 497.345 182.880 ;
    END
  END out1[7]
  PIN out1[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.290 504.065 216.570 508.065 ;
    END
  END out1[8]
  PIN out1[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 504.065 135.610 508.065 ;
    END
  END out1[9]
  PIN out2[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END out2[0]
  PIN out2[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END out2[10]
  PIN out2[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.450 504.065 99.730 508.065 ;
    END
  END out2[11]
  PIN out2[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 137.400 497.345 138.000 ;
    END
  END out2[12]
  PIN out2[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END out2[13]
  PIN out2[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END out2[14]
  PIN out2[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 246.650 504.065 246.930 508.065 ;
    END
  END out2[15]
  PIN out2[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 311.970 504.065 312.250 508.065 ;
    END
  END out2[16]
  PIN out2[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END out2[17]
  PIN out2[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 391.720 497.345 392.320 ;
    END
  END out2[18]
  PIN out2[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END out2[19]
  PIN out2[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END out2[1]
  PIN out2[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.050 504.065 150.330 508.065 ;
    END
  END out2[20]
  PIN out2[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END out2[21]
  PIN out2[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 496.440 497.345 497.040 ;
    END
  END out2[22]
  PIN out2[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END out2[23]
  PIN out2[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 233.960 497.345 234.560 ;
    END
  END out2[24]
  PIN out2[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END out2[25]
  PIN out2[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 47.640 497.345 48.240 ;
    END
  END out2[26]
  PIN out2[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END out2[27]
  PIN out2[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 443.530 504.065 443.810 508.065 ;
    END
  END out2[28]
  PIN out2[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END out2[29]
  PIN out2[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 241.130 504.065 241.410 508.065 ;
    END
  END out2[2]
  PIN out2[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END out2[30]
  PIN out2[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END out2[31]
  PIN out2[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.570 504.065 63.850 508.065 ;
    END
  END out2[3]
  PIN out2[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.930 504.065 393.210 508.065 ;
    END
  END out2[4]
  PIN out2[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.530 504.065 190.810 508.065 ;
    END
  END out2[5]
  PIN out2[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END out2[6]
  PIN out2[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.050 504.065 196.330 508.065 ;
    END
  END out2[7]
  PIN out2[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END out2[8]
  PIN out2[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 62.600 497.345 63.200 ;
    END
  END out2[9]
  PIN out3[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END out3[0]
  PIN out3[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.930 504.065 439.210 508.065 ;
    END
  END out3[10]
  PIN out3[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 281.610 504.065 281.890 508.065 ;
    END
  END out3[11]
  PIN out3[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 352.450 504.065 352.730 508.065 ;
    END
  END out3[12]
  PIN out3[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END out3[13]
  PIN out3[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END out3[14]
  PIN out3[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 287.000 497.345 287.600 ;
    END
  END out3[15]
  PIN out3[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END out3[16]
  PIN out3[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END out3[17]
  PIN out3[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 362.570 504.065 362.850 508.065 ;
    END
  END out3[18]
  PIN out3[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.850 504.065 95.130 508.065 ;
    END
  END out3[19]
  PIN out3[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.970 504.065 59.250 508.065 ;
    END
  END out3[1]
  PIN out3[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END out3[20]
  PIN out3[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END out3[21]
  PIN out3[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END out3[22]
  PIN out3[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 266.890 504.065 267.170 508.065 ;
    END
  END out3[23]
  PIN out3[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END out3[24]
  PIN out3[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 84.360 497.345 84.960 ;
    END
  END out3[25]
  PIN out3[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END out3[26]
  PIN out3[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 504.065 8.650 508.065 ;
    END
  END out3[27]
  PIN out3[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.090 504.065 368.370 508.065 ;
    END
  END out3[28]
  PIN out3[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 408.570 504.065 408.850 508.065 ;
    END
  END out3[29]
  PIN out3[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END out3[2]
  PIN out3[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END out3[30]
  PIN out3[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END out3[31]
  PIN out3[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END out3[3]
  PIN out3[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END out3[4]
  PIN out3[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 231.010 504.065 231.290 508.065 ;
    END
  END out3[5]
  PIN out3[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END out3[6]
  PIN out3[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 493.345 9.560 497.345 10.160 ;
    END
  END out3[7]
  PIN out3[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END out3[8]
  PIN out3[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.530 504.065 489.810 508.065 ;
    END
  END out3[9]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END rst
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 491.740 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 491.740 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 491.740 495.125 ;
      LAYER met1 ;
        RECT 0.070 4.460 494.430 503.840 ;
      LAYER met2 ;
        RECT 0.100 503.785 2.570 504.065 ;
        RECT 3.410 503.785 8.090 504.065 ;
        RECT 8.930 503.785 12.690 504.065 ;
        RECT 13.530 503.785 18.210 504.065 ;
        RECT 19.050 503.785 22.810 504.065 ;
        RECT 23.650 503.785 28.330 504.065 ;
        RECT 29.170 503.785 32.930 504.065 ;
        RECT 33.770 503.785 38.450 504.065 ;
        RECT 39.290 503.785 43.050 504.065 ;
        RECT 43.890 503.785 48.570 504.065 ;
        RECT 49.410 503.785 53.170 504.065 ;
        RECT 54.010 503.785 58.690 504.065 ;
        RECT 59.530 503.785 63.290 504.065 ;
        RECT 64.130 503.785 68.810 504.065 ;
        RECT 69.650 503.785 73.410 504.065 ;
        RECT 74.250 503.785 78.930 504.065 ;
        RECT 79.770 503.785 84.450 504.065 ;
        RECT 85.290 503.785 89.050 504.065 ;
        RECT 89.890 503.785 94.570 504.065 ;
        RECT 95.410 503.785 99.170 504.065 ;
        RECT 100.010 503.785 104.690 504.065 ;
        RECT 105.530 503.785 109.290 504.065 ;
        RECT 110.130 503.785 114.810 504.065 ;
        RECT 115.650 503.785 119.410 504.065 ;
        RECT 120.250 503.785 124.930 504.065 ;
        RECT 125.770 503.785 129.530 504.065 ;
        RECT 130.370 503.785 135.050 504.065 ;
        RECT 135.890 503.785 139.650 504.065 ;
        RECT 140.490 503.785 145.170 504.065 ;
        RECT 146.010 503.785 149.770 504.065 ;
        RECT 150.610 503.785 155.290 504.065 ;
        RECT 156.130 503.785 159.890 504.065 ;
        RECT 160.730 503.785 165.410 504.065 ;
        RECT 166.250 503.785 170.010 504.065 ;
        RECT 170.850 503.785 175.530 504.065 ;
        RECT 176.370 503.785 180.130 504.065 ;
        RECT 180.970 503.785 185.650 504.065 ;
        RECT 186.490 503.785 190.250 504.065 ;
        RECT 191.090 503.785 195.770 504.065 ;
        RECT 196.610 503.785 200.370 504.065 ;
        RECT 201.210 503.785 205.890 504.065 ;
        RECT 206.730 503.785 210.490 504.065 ;
        RECT 211.330 503.785 216.010 504.065 ;
        RECT 216.850 503.785 220.610 504.065 ;
        RECT 221.450 503.785 226.130 504.065 ;
        RECT 226.970 503.785 230.730 504.065 ;
        RECT 231.570 503.785 236.250 504.065 ;
        RECT 237.090 503.785 240.850 504.065 ;
        RECT 241.690 503.785 246.370 504.065 ;
        RECT 247.210 503.785 250.970 504.065 ;
        RECT 251.810 503.785 256.490 504.065 ;
        RECT 257.330 503.785 261.090 504.065 ;
        RECT 261.930 503.785 266.610 504.065 ;
        RECT 267.450 503.785 271.210 504.065 ;
        RECT 272.050 503.785 276.730 504.065 ;
        RECT 277.570 503.785 281.330 504.065 ;
        RECT 282.170 503.785 286.850 504.065 ;
        RECT 287.690 503.785 291.450 504.065 ;
        RECT 292.290 503.785 296.970 504.065 ;
        RECT 297.810 503.785 301.570 504.065 ;
        RECT 302.410 503.785 307.090 504.065 ;
        RECT 307.930 503.785 311.690 504.065 ;
        RECT 312.530 503.785 317.210 504.065 ;
        RECT 318.050 503.785 321.810 504.065 ;
        RECT 322.650 503.785 327.330 504.065 ;
        RECT 328.170 503.785 331.930 504.065 ;
        RECT 332.770 503.785 337.450 504.065 ;
        RECT 338.290 503.785 342.050 504.065 ;
        RECT 342.890 503.785 347.570 504.065 ;
        RECT 348.410 503.785 352.170 504.065 ;
        RECT 353.010 503.785 357.690 504.065 ;
        RECT 358.530 503.785 362.290 504.065 ;
        RECT 363.130 503.785 367.810 504.065 ;
        RECT 368.650 503.785 372.410 504.065 ;
        RECT 373.250 503.785 377.930 504.065 ;
        RECT 378.770 503.785 382.530 504.065 ;
        RECT 383.370 503.785 388.050 504.065 ;
        RECT 388.890 503.785 392.650 504.065 ;
        RECT 393.490 503.785 398.170 504.065 ;
        RECT 399.010 503.785 402.770 504.065 ;
        RECT 403.610 503.785 408.290 504.065 ;
        RECT 409.130 503.785 412.890 504.065 ;
        RECT 413.730 503.785 418.410 504.065 ;
        RECT 419.250 503.785 423.010 504.065 ;
        RECT 423.850 503.785 428.530 504.065 ;
        RECT 429.370 503.785 433.130 504.065 ;
        RECT 433.970 503.785 438.650 504.065 ;
        RECT 439.490 503.785 443.250 504.065 ;
        RECT 444.090 503.785 448.770 504.065 ;
        RECT 449.610 503.785 453.370 504.065 ;
        RECT 454.210 503.785 458.890 504.065 ;
        RECT 459.730 503.785 463.490 504.065 ;
        RECT 464.330 503.785 469.010 504.065 ;
        RECT 469.850 503.785 473.610 504.065 ;
        RECT 474.450 503.785 479.130 504.065 ;
        RECT 479.970 503.785 483.730 504.065 ;
        RECT 484.570 503.785 489.250 504.065 ;
        RECT 490.090 503.785 493.850 504.065 ;
        RECT 0.100 4.280 494.400 503.785 ;
        RECT 0.100 4.000 2.570 4.280 ;
        RECT 3.410 4.000 7.170 4.280 ;
        RECT 8.010 4.000 12.690 4.280 ;
        RECT 13.530 4.000 17.290 4.280 ;
        RECT 18.130 4.000 22.810 4.280 ;
        RECT 23.650 4.000 27.410 4.280 ;
        RECT 28.250 4.000 32.930 4.280 ;
        RECT 33.770 4.000 37.530 4.280 ;
        RECT 38.370 4.000 43.050 4.280 ;
        RECT 43.890 4.000 47.650 4.280 ;
        RECT 48.490 4.000 53.170 4.280 ;
        RECT 54.010 4.000 57.770 4.280 ;
        RECT 58.610 4.000 63.290 4.280 ;
        RECT 64.130 4.000 67.890 4.280 ;
        RECT 68.730 4.000 73.410 4.280 ;
        RECT 74.250 4.000 78.010 4.280 ;
        RECT 78.850 4.000 83.530 4.280 ;
        RECT 84.370 4.000 88.130 4.280 ;
        RECT 88.970 4.000 93.650 4.280 ;
        RECT 94.490 4.000 98.250 4.280 ;
        RECT 99.090 4.000 103.770 4.280 ;
        RECT 104.610 4.000 108.370 4.280 ;
        RECT 109.210 4.000 113.890 4.280 ;
        RECT 114.730 4.000 118.490 4.280 ;
        RECT 119.330 4.000 124.010 4.280 ;
        RECT 124.850 4.000 128.610 4.280 ;
        RECT 129.450 4.000 134.130 4.280 ;
        RECT 134.970 4.000 138.730 4.280 ;
        RECT 139.570 4.000 144.250 4.280 ;
        RECT 145.090 4.000 148.850 4.280 ;
        RECT 149.690 4.000 154.370 4.280 ;
        RECT 155.210 4.000 158.970 4.280 ;
        RECT 159.810 4.000 164.490 4.280 ;
        RECT 165.330 4.000 169.090 4.280 ;
        RECT 169.930 4.000 174.610 4.280 ;
        RECT 175.450 4.000 179.210 4.280 ;
        RECT 180.050 4.000 184.730 4.280 ;
        RECT 185.570 4.000 189.330 4.280 ;
        RECT 190.170 4.000 194.850 4.280 ;
        RECT 195.690 4.000 199.450 4.280 ;
        RECT 200.290 4.000 204.970 4.280 ;
        RECT 205.810 4.000 209.570 4.280 ;
        RECT 210.410 4.000 215.090 4.280 ;
        RECT 215.930 4.000 219.690 4.280 ;
        RECT 220.530 4.000 225.210 4.280 ;
        RECT 226.050 4.000 229.810 4.280 ;
        RECT 230.650 4.000 235.330 4.280 ;
        RECT 236.170 4.000 239.930 4.280 ;
        RECT 240.770 4.000 245.450 4.280 ;
        RECT 246.290 4.000 250.050 4.280 ;
        RECT 250.890 4.000 255.570 4.280 ;
        RECT 256.410 4.000 260.170 4.280 ;
        RECT 261.010 4.000 265.690 4.280 ;
        RECT 266.530 4.000 270.290 4.280 ;
        RECT 271.130 4.000 275.810 4.280 ;
        RECT 276.650 4.000 280.410 4.280 ;
        RECT 281.250 4.000 285.930 4.280 ;
        RECT 286.770 4.000 290.530 4.280 ;
        RECT 291.370 4.000 296.050 4.280 ;
        RECT 296.890 4.000 300.650 4.280 ;
        RECT 301.490 4.000 306.170 4.280 ;
        RECT 307.010 4.000 310.770 4.280 ;
        RECT 311.610 4.000 316.290 4.280 ;
        RECT 317.130 4.000 320.890 4.280 ;
        RECT 321.730 4.000 326.410 4.280 ;
        RECT 327.250 4.000 331.010 4.280 ;
        RECT 331.850 4.000 336.530 4.280 ;
        RECT 337.370 4.000 341.130 4.280 ;
        RECT 341.970 4.000 346.650 4.280 ;
        RECT 347.490 4.000 351.250 4.280 ;
        RECT 352.090 4.000 356.770 4.280 ;
        RECT 357.610 4.000 361.370 4.280 ;
        RECT 362.210 4.000 366.890 4.280 ;
        RECT 367.730 4.000 371.490 4.280 ;
        RECT 372.330 4.000 377.010 4.280 ;
        RECT 377.850 4.000 381.610 4.280 ;
        RECT 382.450 4.000 387.130 4.280 ;
        RECT 387.970 4.000 391.730 4.280 ;
        RECT 392.570 4.000 397.250 4.280 ;
        RECT 398.090 4.000 401.850 4.280 ;
        RECT 402.690 4.000 407.370 4.280 ;
        RECT 408.210 4.000 411.970 4.280 ;
        RECT 412.810 4.000 417.490 4.280 ;
        RECT 418.330 4.000 423.010 4.280 ;
        RECT 423.850 4.000 427.610 4.280 ;
        RECT 428.450 4.000 433.130 4.280 ;
        RECT 433.970 4.000 437.730 4.280 ;
        RECT 438.570 4.000 443.250 4.280 ;
        RECT 444.090 4.000 447.850 4.280 ;
        RECT 448.690 4.000 453.370 4.280 ;
        RECT 454.210 4.000 457.970 4.280 ;
        RECT 458.810 4.000 463.490 4.280 ;
        RECT 464.330 4.000 468.090 4.280 ;
        RECT 468.930 4.000 473.610 4.280 ;
        RECT 474.450 4.000 478.210 4.280 ;
        RECT 479.050 4.000 483.730 4.280 ;
        RECT 484.570 4.000 488.330 4.280 ;
        RECT 489.170 4.000 493.850 4.280 ;
      LAYER met3 ;
        RECT 4.400 497.440 493.345 498.265 ;
        RECT 4.400 497.400 492.945 497.440 ;
        RECT 3.990 496.040 492.945 497.400 ;
        RECT 3.990 490.640 493.345 496.040 ;
        RECT 4.400 489.280 493.345 490.640 ;
        RECT 4.400 489.240 492.945 489.280 ;
        RECT 3.990 487.880 492.945 489.240 ;
        RECT 3.990 483.840 493.345 487.880 ;
        RECT 4.400 482.480 493.345 483.840 ;
        RECT 4.400 482.440 492.945 482.480 ;
        RECT 3.990 481.080 492.945 482.440 ;
        RECT 3.990 475.680 493.345 481.080 ;
        RECT 4.400 474.320 493.345 475.680 ;
        RECT 4.400 474.280 492.945 474.320 ;
        RECT 3.990 472.920 492.945 474.280 ;
        RECT 3.990 468.880 493.345 472.920 ;
        RECT 4.400 467.520 493.345 468.880 ;
        RECT 4.400 467.480 492.945 467.520 ;
        RECT 3.990 466.120 492.945 467.480 ;
        RECT 3.990 460.720 493.345 466.120 ;
        RECT 4.400 459.360 493.345 460.720 ;
        RECT 4.400 459.320 492.945 459.360 ;
        RECT 3.990 457.960 492.945 459.320 ;
        RECT 3.990 453.920 493.345 457.960 ;
        RECT 4.400 452.560 493.345 453.920 ;
        RECT 4.400 452.520 492.945 452.560 ;
        RECT 3.990 451.160 492.945 452.520 ;
        RECT 3.990 445.760 493.345 451.160 ;
        RECT 4.400 444.400 493.345 445.760 ;
        RECT 4.400 444.360 492.945 444.400 ;
        RECT 3.990 443.000 492.945 444.360 ;
        RECT 3.990 438.960 493.345 443.000 ;
        RECT 4.400 437.600 493.345 438.960 ;
        RECT 4.400 437.560 492.945 437.600 ;
        RECT 3.990 436.200 492.945 437.560 ;
        RECT 3.990 430.800 493.345 436.200 ;
        RECT 4.400 429.440 493.345 430.800 ;
        RECT 4.400 429.400 492.945 429.440 ;
        RECT 3.990 428.040 492.945 429.400 ;
        RECT 3.990 424.000 493.345 428.040 ;
        RECT 4.400 422.640 493.345 424.000 ;
        RECT 4.400 422.600 492.945 422.640 ;
        RECT 3.990 421.240 492.945 422.600 ;
        RECT 3.990 415.840 493.345 421.240 ;
        RECT 4.400 414.480 493.345 415.840 ;
        RECT 4.400 414.440 492.945 414.480 ;
        RECT 3.990 413.080 492.945 414.440 ;
        RECT 3.990 409.040 493.345 413.080 ;
        RECT 4.400 407.680 493.345 409.040 ;
        RECT 4.400 407.640 492.945 407.680 ;
        RECT 3.990 406.280 492.945 407.640 ;
        RECT 3.990 400.880 493.345 406.280 ;
        RECT 4.400 399.520 493.345 400.880 ;
        RECT 4.400 399.480 492.945 399.520 ;
        RECT 3.990 398.120 492.945 399.480 ;
        RECT 3.990 394.080 493.345 398.120 ;
        RECT 4.400 392.720 493.345 394.080 ;
        RECT 4.400 392.680 492.945 392.720 ;
        RECT 3.990 391.320 492.945 392.680 ;
        RECT 3.990 385.920 493.345 391.320 ;
        RECT 4.400 384.560 493.345 385.920 ;
        RECT 4.400 384.520 492.945 384.560 ;
        RECT 3.990 383.160 492.945 384.520 ;
        RECT 3.990 379.120 493.345 383.160 ;
        RECT 4.400 377.760 493.345 379.120 ;
        RECT 4.400 377.720 492.945 377.760 ;
        RECT 3.990 376.360 492.945 377.720 ;
        RECT 3.990 370.960 493.345 376.360 ;
        RECT 4.400 369.600 493.345 370.960 ;
        RECT 4.400 369.560 492.945 369.600 ;
        RECT 3.990 368.200 492.945 369.560 ;
        RECT 3.990 364.160 493.345 368.200 ;
        RECT 4.400 362.800 493.345 364.160 ;
        RECT 4.400 362.760 492.945 362.800 ;
        RECT 3.990 361.400 492.945 362.760 ;
        RECT 3.990 356.000 493.345 361.400 ;
        RECT 4.400 354.640 493.345 356.000 ;
        RECT 4.400 354.600 492.945 354.640 ;
        RECT 3.990 353.240 492.945 354.600 ;
        RECT 3.990 349.200 493.345 353.240 ;
        RECT 4.400 347.840 493.345 349.200 ;
        RECT 4.400 347.800 492.945 347.840 ;
        RECT 3.990 346.440 492.945 347.800 ;
        RECT 3.990 341.040 493.345 346.440 ;
        RECT 4.400 339.680 493.345 341.040 ;
        RECT 4.400 339.640 492.945 339.680 ;
        RECT 3.990 338.280 492.945 339.640 ;
        RECT 3.990 334.240 493.345 338.280 ;
        RECT 4.400 332.880 493.345 334.240 ;
        RECT 4.400 332.840 492.945 332.880 ;
        RECT 3.990 331.480 492.945 332.840 ;
        RECT 3.990 326.080 493.345 331.480 ;
        RECT 4.400 324.720 493.345 326.080 ;
        RECT 4.400 324.680 492.945 324.720 ;
        RECT 3.990 323.320 492.945 324.680 ;
        RECT 3.990 319.280 493.345 323.320 ;
        RECT 4.400 317.920 493.345 319.280 ;
        RECT 4.400 317.880 492.945 317.920 ;
        RECT 3.990 316.520 492.945 317.880 ;
        RECT 3.990 311.120 493.345 316.520 ;
        RECT 4.400 309.760 493.345 311.120 ;
        RECT 4.400 309.720 492.945 309.760 ;
        RECT 3.990 308.360 492.945 309.720 ;
        RECT 3.990 304.320 493.345 308.360 ;
        RECT 4.400 302.960 493.345 304.320 ;
        RECT 4.400 302.920 492.945 302.960 ;
        RECT 3.990 301.560 492.945 302.920 ;
        RECT 3.990 296.160 493.345 301.560 ;
        RECT 4.400 294.800 493.345 296.160 ;
        RECT 4.400 294.760 492.945 294.800 ;
        RECT 3.990 293.400 492.945 294.760 ;
        RECT 3.990 289.360 493.345 293.400 ;
        RECT 4.400 288.000 493.345 289.360 ;
        RECT 4.400 287.960 492.945 288.000 ;
        RECT 3.990 286.600 492.945 287.960 ;
        RECT 3.990 281.200 493.345 286.600 ;
        RECT 4.400 279.840 493.345 281.200 ;
        RECT 4.400 279.800 492.945 279.840 ;
        RECT 3.990 278.440 492.945 279.800 ;
        RECT 3.990 274.400 493.345 278.440 ;
        RECT 4.400 273.040 493.345 274.400 ;
        RECT 4.400 273.000 492.945 273.040 ;
        RECT 3.990 271.640 492.945 273.000 ;
        RECT 3.990 266.240 493.345 271.640 ;
        RECT 4.400 264.880 493.345 266.240 ;
        RECT 4.400 264.840 492.945 264.880 ;
        RECT 3.990 263.480 492.945 264.840 ;
        RECT 3.990 259.440 493.345 263.480 ;
        RECT 4.400 258.080 493.345 259.440 ;
        RECT 4.400 258.040 492.945 258.080 ;
        RECT 3.990 256.680 492.945 258.040 ;
        RECT 3.990 251.280 493.345 256.680 ;
        RECT 4.400 249.920 493.345 251.280 ;
        RECT 4.400 249.880 492.945 249.920 ;
        RECT 3.990 248.520 492.945 249.880 ;
        RECT 3.990 244.480 493.345 248.520 ;
        RECT 4.400 243.120 493.345 244.480 ;
        RECT 4.400 243.080 492.945 243.120 ;
        RECT 3.990 241.720 492.945 243.080 ;
        RECT 3.990 236.320 493.345 241.720 ;
        RECT 4.400 234.960 493.345 236.320 ;
        RECT 4.400 234.920 492.945 234.960 ;
        RECT 3.990 233.560 492.945 234.920 ;
        RECT 3.990 229.520 493.345 233.560 ;
        RECT 4.400 228.160 493.345 229.520 ;
        RECT 4.400 228.120 492.945 228.160 ;
        RECT 3.990 226.760 492.945 228.120 ;
        RECT 3.990 221.360 493.345 226.760 ;
        RECT 4.400 220.000 493.345 221.360 ;
        RECT 4.400 219.960 492.945 220.000 ;
        RECT 3.990 218.600 492.945 219.960 ;
        RECT 3.990 214.560 493.345 218.600 ;
        RECT 4.400 213.200 493.345 214.560 ;
        RECT 4.400 213.160 492.945 213.200 ;
        RECT 3.990 211.800 492.945 213.160 ;
        RECT 3.990 206.400 493.345 211.800 ;
        RECT 4.400 205.040 493.345 206.400 ;
        RECT 4.400 205.000 492.945 205.040 ;
        RECT 3.990 203.640 492.945 205.000 ;
        RECT 3.990 199.600 493.345 203.640 ;
        RECT 4.400 198.240 493.345 199.600 ;
        RECT 4.400 198.200 492.945 198.240 ;
        RECT 3.990 196.840 492.945 198.200 ;
        RECT 3.990 191.440 493.345 196.840 ;
        RECT 4.400 190.080 493.345 191.440 ;
        RECT 4.400 190.040 492.945 190.080 ;
        RECT 3.990 188.680 492.945 190.040 ;
        RECT 3.990 184.640 493.345 188.680 ;
        RECT 4.400 183.280 493.345 184.640 ;
        RECT 4.400 183.240 492.945 183.280 ;
        RECT 3.990 181.880 492.945 183.240 ;
        RECT 3.990 176.480 493.345 181.880 ;
        RECT 4.400 175.120 493.345 176.480 ;
        RECT 4.400 175.080 492.945 175.120 ;
        RECT 3.990 173.720 492.945 175.080 ;
        RECT 3.990 169.680 493.345 173.720 ;
        RECT 4.400 168.320 493.345 169.680 ;
        RECT 4.400 168.280 492.945 168.320 ;
        RECT 3.990 166.920 492.945 168.280 ;
        RECT 3.990 161.520 493.345 166.920 ;
        RECT 4.400 160.160 493.345 161.520 ;
        RECT 4.400 160.120 492.945 160.160 ;
        RECT 3.990 158.760 492.945 160.120 ;
        RECT 3.990 154.720 493.345 158.760 ;
        RECT 4.400 153.360 493.345 154.720 ;
        RECT 4.400 153.320 492.945 153.360 ;
        RECT 3.990 151.960 492.945 153.320 ;
        RECT 3.990 146.560 493.345 151.960 ;
        RECT 4.400 145.200 493.345 146.560 ;
        RECT 4.400 145.160 492.945 145.200 ;
        RECT 3.990 143.800 492.945 145.160 ;
        RECT 3.990 139.760 493.345 143.800 ;
        RECT 4.400 138.400 493.345 139.760 ;
        RECT 4.400 138.360 492.945 138.400 ;
        RECT 3.990 137.000 492.945 138.360 ;
        RECT 3.990 131.600 493.345 137.000 ;
        RECT 4.400 130.240 493.345 131.600 ;
        RECT 4.400 130.200 492.945 130.240 ;
        RECT 3.990 128.840 492.945 130.200 ;
        RECT 3.990 124.800 493.345 128.840 ;
        RECT 4.400 123.440 493.345 124.800 ;
        RECT 4.400 123.400 492.945 123.440 ;
        RECT 3.990 122.040 492.945 123.400 ;
        RECT 3.990 116.640 493.345 122.040 ;
        RECT 4.400 115.280 493.345 116.640 ;
        RECT 4.400 115.240 492.945 115.280 ;
        RECT 3.990 113.880 492.945 115.240 ;
        RECT 3.990 109.840 493.345 113.880 ;
        RECT 4.400 108.480 493.345 109.840 ;
        RECT 4.400 108.440 492.945 108.480 ;
        RECT 3.990 107.080 492.945 108.440 ;
        RECT 3.990 101.680 493.345 107.080 ;
        RECT 4.400 100.320 493.345 101.680 ;
        RECT 4.400 100.280 492.945 100.320 ;
        RECT 3.990 98.920 492.945 100.280 ;
        RECT 3.990 94.880 493.345 98.920 ;
        RECT 4.400 93.520 493.345 94.880 ;
        RECT 4.400 93.480 492.945 93.520 ;
        RECT 3.990 92.120 492.945 93.480 ;
        RECT 3.990 86.720 493.345 92.120 ;
        RECT 4.400 85.360 493.345 86.720 ;
        RECT 4.400 85.320 492.945 85.360 ;
        RECT 3.990 83.960 492.945 85.320 ;
        RECT 3.990 79.920 493.345 83.960 ;
        RECT 4.400 78.560 493.345 79.920 ;
        RECT 4.400 78.520 492.945 78.560 ;
        RECT 3.990 77.160 492.945 78.520 ;
        RECT 3.990 71.760 493.345 77.160 ;
        RECT 4.400 70.400 493.345 71.760 ;
        RECT 4.400 70.360 492.945 70.400 ;
        RECT 3.990 69.000 492.945 70.360 ;
        RECT 3.990 64.960 493.345 69.000 ;
        RECT 4.400 63.600 493.345 64.960 ;
        RECT 4.400 63.560 492.945 63.600 ;
        RECT 3.990 62.200 492.945 63.560 ;
        RECT 3.990 56.800 493.345 62.200 ;
        RECT 4.400 55.440 493.345 56.800 ;
        RECT 4.400 55.400 492.945 55.440 ;
        RECT 3.990 54.040 492.945 55.400 ;
        RECT 3.990 50.000 493.345 54.040 ;
        RECT 4.400 48.640 493.345 50.000 ;
        RECT 4.400 48.600 492.945 48.640 ;
        RECT 3.990 47.240 492.945 48.600 ;
        RECT 3.990 41.840 493.345 47.240 ;
        RECT 4.400 40.480 493.345 41.840 ;
        RECT 4.400 40.440 492.945 40.480 ;
        RECT 3.990 39.080 492.945 40.440 ;
        RECT 3.990 35.040 493.345 39.080 ;
        RECT 4.400 33.680 493.345 35.040 ;
        RECT 4.400 33.640 492.945 33.680 ;
        RECT 3.990 32.280 492.945 33.640 ;
        RECT 3.990 26.880 493.345 32.280 ;
        RECT 4.400 25.520 493.345 26.880 ;
        RECT 4.400 25.480 492.945 25.520 ;
        RECT 3.990 24.120 492.945 25.480 ;
        RECT 3.990 20.080 493.345 24.120 ;
        RECT 4.400 18.720 493.345 20.080 ;
        RECT 4.400 18.680 492.945 18.720 ;
        RECT 3.990 17.320 492.945 18.680 ;
        RECT 3.990 11.920 493.345 17.320 ;
        RECT 4.400 10.560 493.345 11.920 ;
        RECT 4.400 10.520 492.945 10.560 ;
        RECT 3.990 9.160 492.945 10.520 ;
        RECT 3.990 4.255 493.345 9.160 ;
      LAYER met4 ;
        RECT 11.335 10.640 483.440 495.280 ;
      LAYER met5 ;
        RECT 5.520 179.670 491.740 487.630 ;
  END
END mac_cluster
END LIBRARY

