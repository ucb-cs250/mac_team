`define SINGLE 0
`define DUAL 1
`define QUAD 2