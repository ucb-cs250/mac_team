VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mac_cluster
  CLASS BLOCK ;
  FOREIGN mac_cluster ;
  ORIGIN 0.000 0.000 ;
  SIZE 479.500 BY 490.220 ;
  PIN A0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.570 486.220 178.850 490.220 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 261.160 479.500 261.760 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.050 486.220 403.330 490.220 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.290 486.220 193.570 490.220 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END A0[7]
  PIN A1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.370 486.220 169.650 490.220 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 448.840 479.500 449.440 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 252.170 486.220 252.450 490.220 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 276.090 486.220 276.370 490.220 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 486.220 17.850 490.220 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 261.370 486.220 261.650 490.220 ;
    END
  END A1[7]
  PIN A2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.490 486.220 432.770 490.220 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END A2[6]
  PIN A2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 427.080 479.500 427.680 ;
    END
  END A2[7]
  PIN A3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.330 486.220 227.610 490.220 ;
    END
  END A3[0]
  PIN A3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END A3[1]
  PIN A3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 447.210 486.220 447.490 490.220 ;
    END
  END A3[2]
  PIN A3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 197.890 486.220 198.170 490.220 ;
    END
  END A3[3]
  PIN A3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END A3[4]
  PIN A3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END A3[5]
  PIN A3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END A3[6]
  PIN A3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.330 486.220 66.610 490.220 ;
    END
  END A3[7]
  PIN B0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END B0[0]
  PIN B0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END B0[1]
  PIN B0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END B0[2]
  PIN B0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END B0[3]
  PIN B0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 210.840 479.500 211.440 ;
    END
  END B0[4]
  PIN B0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.130 486.220 218.410 490.220 ;
    END
  END B0[5]
  PIN B0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 486.220 72.130 490.220 ;
    END
  END B0[6]
  PIN B0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END B0[7]
  PIN B1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.930 486.220 140.210 490.220 ;
    END
  END B1[0]
  PIN B1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 355.000 479.500 355.600 ;
    END
  END B1[1]
  PIN B1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 145.560 479.500 146.160 ;
    END
  END B1[2]
  PIN B1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END B1[3]
  PIN B1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 358.890 486.220 359.170 490.220 ;
    END
  END B1[4]
  PIN B1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END B1[5]
  PIN B1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.130 486.220 149.410 490.220 ;
    END
  END B1[6]
  PIN B1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 232.600 479.500 233.200 ;
    END
  END B1[7]
  PIN B2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END B2[0]
  PIN B2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END B2[1]
  PIN B2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END B2[2]
  PIN B2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 110.200 479.500 110.800 ;
    END
  END B2[3]
  PIN B2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.650 486.220 154.930 490.220 ;
    END
  END B2[4]
  PIN B2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 486.220 23.370 490.220 ;
    END
  END B2[5]
  PIN B2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END B2[6]
  PIN B2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 269.320 479.500 269.920 ;
    END
  END B2[7]
  PIN B3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 73.480 479.500 74.080 ;
    END
  END B3[0]
  PIN B3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END B3[1]
  PIN B3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END B3[2]
  PIN B3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 463.800 479.500 464.400 ;
    END
  END B3[3]
  PIN B3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 204.040 479.500 204.640 ;
    END
  END B3[4]
  PIN B3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.690 486.220 27.970 490.220 ;
    END
  END B3[5]
  PIN B3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END B3[6]
  PIN B3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 103.400 479.500 104.000 ;
    END
  END B3[7]
  PIN cfg[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.650 486.220 246.930 490.220 ;
    END
  END cfg[0]
  PIN cfg[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END cfg[100]
  PIN cfg[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END cfg[101]
  PIN cfg[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END cfg[102]
  PIN cfg[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 486.220 47.290 490.220 ;
    END
  END cfg[103]
  PIN cfg[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END cfg[104]
  PIN cfg[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END cfg[105]
  PIN cfg[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 413.480 479.500 414.080 ;
    END
  END cfg[106]
  PIN cfg[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END cfg[107]
  PIN cfg[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END cfg[108]
  PIN cfg[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 486.220 106.170 490.220 ;
    END
  END cfg[109]
  PIN cfg[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END cfg[10]
  PIN cfg[110]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END cfg[110]
  PIN cfg[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END cfg[111]
  PIN cfg[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END cfg[112]
  PIN cfg[113]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 197.240 479.500 197.840 ;
    END
  END cfg[113]
  PIN cfg[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 239.400 479.500 240.000 ;
    END
  END cfg[114]
  PIN cfg[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.570 486.220 86.850 490.220 ;
    END
  END cfg[115]
  PIN cfg[116]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END cfg[116]
  PIN cfg[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 413.170 486.220 413.450 490.220 ;
    END
  END cfg[117]
  PIN cfg[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END cfg[118]
  PIN cfg[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END cfg[119]
  PIN cfg[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END cfg[11]
  PIN cfg[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 486.220 115.370 490.220 ;
    END
  END cfg[120]
  PIN cfg[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 23.160 479.500 23.760 ;
    END
  END cfg[121]
  PIN cfg[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END cfg[122]
  PIN cfg[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END cfg[123]
  PIN cfg[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 348.200 479.500 348.800 ;
    END
  END cfg[124]
  PIN cfg[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 486.220 32.570 490.220 ;
    END
  END cfg[125]
  PIN cfg[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 247.560 479.500 248.160 ;
    END
  END cfg[126]
  PIN cfg[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END cfg[127]
  PIN cfg[128]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END cfg[128]
  PIN cfg[129]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END cfg[129]
  PIN cfg[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END cfg[12]
  PIN cfg[130]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END cfg[130]
  PIN cfg[131]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.970 486.220 335.250 490.220 ;
    END
  END cfg[131]
  PIN cfg[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 310.130 486.220 310.410 490.220 ;
    END
  END cfg[13]
  PIN cfg[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END cfg[14]
  PIN cfg[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END cfg[15]
  PIN cfg[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END cfg[16]
  PIN cfg[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.610 486.220 281.890 490.220 ;
    END
  END cfg[17]
  PIN cfg[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 341.400 479.500 342.000 ;
    END
  END cfg[18]
  PIN cfg[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END cfg[19]
  PIN cfg[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END cfg[1]
  PIN cfg[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 203.410 486.220 203.690 490.220 ;
    END
  END cfg[20]
  PIN cfg[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 88.440 479.500 89.040 ;
    END
  END cfg[21]
  PIN cfg[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 167.320 479.500 167.920 ;
    END
  END cfg[22]
  PIN cfg[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END cfg[23]
  PIN cfg[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 16.360 479.500 16.960 ;
    END
  END cfg[24]
  PIN cfg[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END cfg[25]
  PIN cfg[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END cfg[26]
  PIN cfg[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 324.850 486.220 325.130 490.220 ;
    END
  END cfg[27]
  PIN cfg[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 417.770 486.220 418.050 490.220 ;
    END
  END cfg[28]
  PIN cfg[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END cfg[29]
  PIN cfg[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END cfg[2]
  PIN cfg[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END cfg[30]
  PIN cfg[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 304.680 479.500 305.280 ;
    END
  END cfg[31]
  PIN cfg[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 451.810 486.220 452.090 490.220 ;
    END
  END cfg[32]
  PIN cfg[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.050 486.220 242.330 490.220 ;
    END
  END cfg[33]
  PIN cfg[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END cfg[34]
  PIN cfg[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END cfg[35]
  PIN cfg[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END cfg[36]
  PIN cfg[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END cfg[37]
  PIN cfg[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 53.080 479.500 53.680 ;
    END
  END cfg[38]
  PIN cfg[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 369.960 479.500 370.560 ;
    END
  END cfg[39]
  PIN cfg[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 442.040 479.500 442.640 ;
    END
  END cfg[3]
  PIN cfg[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END cfg[40]
  PIN cfg[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.050 486.220 81.330 490.220 ;
    END
  END cfg[41]
  PIN cfg[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END cfg[42]
  PIN cfg[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END cfg[43]
  PIN cfg[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 125.160 479.500 125.760 ;
    END
  END cfg[44]
  PIN cfg[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END cfg[45]
  PIN cfg[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 391.720 479.500 392.320 ;
    END
  END cfg[46]
  PIN cfg[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.730 486.220 384.010 490.220 ;
    END
  END cfg[47]
  PIN cfg[48]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END cfg[48]
  PIN cfg[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.450 486.220 76.730 490.220 ;
    END
  END cfg[49]
  PIN cfg[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 163.850 486.220 164.130 490.220 ;
    END
  END cfg[4]
  PIN cfg[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END cfg[50]
  PIN cfg[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 441.690 486.220 441.970 490.220 ;
    END
  END cfg[51]
  PIN cfg[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END cfg[52]
  PIN cfg[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END cfg[53]
  PIN cfg[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END cfg[54]
  PIN cfg[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END cfg[55]
  PIN cfg[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END cfg[56]
  PIN cfg[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END cfg[57]
  PIN cfg[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 369.010 486.220 369.290 490.220 ;
    END
  END cfg[58]
  PIN cfg[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END cfg[59]
  PIN cfg[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 373.610 486.220 373.890 490.220 ;
    END
  END cfg[5]
  PIN cfg[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 470.600 479.500 471.200 ;
    END
  END cfg[60]
  PIN cfg[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 282.920 479.500 283.520 ;
    END
  END cfg[61]
  PIN cfg[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 286.210 486.220 286.490 490.220 ;
    END
  END cfg[62]
  PIN cfg[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 138.760 479.500 139.360 ;
    END
  END cfg[63]
  PIN cfg[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END cfg[64]
  PIN cfg[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END cfg[65]
  PIN cfg[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 486.220 100.650 490.220 ;
    END
  END cfg[66]
  PIN cfg[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 486.220 4.050 490.220 ;
    END
  END cfg[67]
  PIN cfg[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END cfg[68]
  PIN cfg[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END cfg[69]
  PIN cfg[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 290.810 486.220 291.090 490.220 ;
    END
  END cfg[6]
  PIN cfg[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END cfg[70]
  PIN cfg[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 153.720 479.500 154.320 ;
    END
  END cfg[71]
  PIN cfg[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END cfg[72]
  PIN cfg[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END cfg[73]
  PIN cfg[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.250 486.220 159.530 490.220 ;
    END
  END cfg[74]
  PIN cfg[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END cfg[75]
  PIN cfg[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END cfg[76]
  PIN cfg[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END cfg[77]
  PIN cfg[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 31.320 479.500 31.920 ;
    END
  END cfg[78]
  PIN cfg[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 388.330 486.220 388.610 490.220 ;
    END
  END cfg[79]
  PIN cfg[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END cfg[7]
  PIN cfg[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END cfg[80]
  PIN cfg[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END cfg[81]
  PIN cfg[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END cfg[82]
  PIN cfg[83]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END cfg[83]
  PIN cfg[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 475.730 486.220 476.010 490.220 ;
    END
  END cfg[84]
  PIN cfg[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 344.170 486.220 344.450 490.220 ;
    END
  END cfg[85]
  PIN cfg[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 305.530 486.220 305.810 490.220 ;
    END
  END cfg[86]
  PIN cfg[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 189.080 479.500 189.680 ;
    END
  END cfg[87]
  PIN cfg[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 320.250 486.220 320.530 490.220 ;
    END
  END cfg[88]
  PIN cfg[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END cfg[89]
  PIN cfg[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 319.640 479.500 320.240 ;
    END
  END cfg[8]
  PIN cfg[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END cfg[90]
  PIN cfg[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END cfg[91]
  PIN cfg[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END cfg[92]
  PIN cfg[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END cfg[93]
  PIN cfg[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END cfg[94]
  PIN cfg[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 486.220 110.770 490.220 ;
    END
  END cfg[95]
  PIN cfg[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 95.240 479.500 95.840 ;
    END
  END cfg[96]
  PIN cfg[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END cfg[97]
  PIN cfg[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END cfg[98]
  PIN cfg[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END cfg[99]
  PIN cfg[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 398.520 479.500 399.120 ;
    END
  END cfg[9]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 456.410 486.220 456.690 490.220 ;
    END
  END clk
  PIN cset
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.500 217.640 479.500 218.240 ;
    END
  END cset
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 266.890 486.220 267.170 490.220 ;
    END
  END en
  PIN out0[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END out0[0]
  PIN out0[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 398.450 486.220 398.730 490.220 ;
    END
  END out0[10]
  PIN out0[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 254.360 479.500 254.960 ;
    END
  END out0[11]
  PIN out0[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 405.320 479.500 405.920 ;
    END
  END out0[12]
  PIN out0[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 289.720 479.500 290.320 ;
    END
  END out0[13]
  PIN out0[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 117.000 479.500 117.600 ;
    END
  END out0[14]
  PIN out0[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 173.970 486.220 174.250 490.220 ;
    END
  END out0[15]
  PIN out0[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 486.220 135.610 490.220 ;
    END
  END out0[16]
  PIN out0[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 486.220 120.890 490.220 ;
    END
  END out0[17]
  PIN out0[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END out0[18]
  PIN out0[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END out0[19]
  PIN out0[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 326.440 479.500 327.040 ;
    END
  END out0[1]
  PIN out0[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END out0[20]
  PIN out0[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END out0[21]
  PIN out0[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END out0[22]
  PIN out0[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END out0[23]
  PIN out0[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.610 486.220 212.890 490.220 ;
    END
  END out0[24]
  PIN out0[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.410 486.220 364.690 490.220 ;
    END
  END out0[25]
  PIN out0[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 383.560 479.500 384.160 ;
    END
  END out0[26]
  PIN out0[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 433.880 479.500 434.480 ;
    END
  END out0[27]
  PIN out0[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.530 486.220 52.810 490.220 ;
    END
  END out0[28]
  PIN out0[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 311.480 479.500 312.080 ;
    END
  END out0[29]
  PIN out0[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 437.090 486.220 437.370 490.220 ;
    END
  END out0[2]
  PIN out0[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END out0[30]
  PIN out0[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END out0[31]
  PIN out0[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END out0[3]
  PIN out0[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 38.120 479.500 38.720 ;
    END
  END out0[4]
  PIN out0[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 361.800 479.500 362.400 ;
    END
  END out0[5]
  PIN out0[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 330.370 486.220 330.650 490.220 ;
    END
  END out0[6]
  PIN out0[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 297.880 479.500 298.480 ;
    END
  END out0[7]
  PIN out0[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END out0[8]
  PIN out0[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.530 486.220 466.810 490.220 ;
    END
  END out0[9]
  PIN out1[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 315.650 486.220 315.930 490.220 ;
    END
  END out1[0]
  PIN out1[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 333.240 479.500 333.840 ;
    END
  END out1[10]
  PIN out1[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 420.280 479.500 420.880 ;
    END
  END out1[11]
  PIN out1[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END out1[12]
  PIN out1[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END out1[13]
  PIN out1[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.410 486.220 42.690 490.220 ;
    END
  END out1[14]
  PIN out1[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.410 486.220 295.690 490.220 ;
    END
  END out1[15]
  PIN out1[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END out1[16]
  PIN out1[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 182.280 479.500 182.880 ;
    END
  END out1[17]
  PIN out1[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 486.220 38.090 490.220 ;
    END
  END out1[18]
  PIN out1[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END out1[19]
  PIN out1[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END out1[1]
  PIN out1[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 455.640 479.500 456.240 ;
    END
  END out1[20]
  PIN out1[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 407.650 486.220 407.930 490.220 ;
    END
  END out1[21]
  PIN out1[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END out1[22]
  PIN out1[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END out1[23]
  PIN out1[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 125.210 486.220 125.490 490.220 ;
    END
  END out1[24]
  PIN out1[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END out1[25]
  PIN out1[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END out1[26]
  PIN out1[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 461.930 486.220 462.210 490.220 ;
    END
  END out1[27]
  PIN out1[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 160.520 479.500 161.120 ;
    END
  END out1[28]
  PIN out1[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END out1[29]
  PIN out1[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END out1[2]
  PIN out1[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END out1[30]
  PIN out1[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.970 486.220 13.250 490.220 ;
    END
  END out1[31]
  PIN out1[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 66.680 479.500 67.280 ;
    END
  END out1[3]
  PIN out1[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END out1[4]
  PIN out1[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END out1[5]
  PIN out1[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END out1[6]
  PIN out1[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 175.480 479.500 176.080 ;
    END
  END out1[7]
  PIN out1[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.010 486.220 208.290 490.220 ;
    END
  END out1[8]
  PIN out1[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 486.220 130.090 490.220 ;
    END
  END out1[9]
  PIN out2[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END out2[0]
  PIN out2[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END out2[10]
  PIN out2[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 486.220 96.050 490.220 ;
    END
  END out2[11]
  PIN out2[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 131.960 479.500 132.560 ;
    END
  END out2[12]
  PIN out2[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END out2[13]
  PIN out2[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END out2[14]
  PIN out2[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 237.450 486.220 237.730 490.220 ;
    END
  END out2[15]
  PIN out2[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 300.930 486.220 301.210 490.220 ;
    END
  END out2[16]
  PIN out2[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END out2[17]
  PIN out2[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 376.760 479.500 377.360 ;
    END
  END out2[18]
  PIN out2[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END out2[19]
  PIN out2[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END out2[1]
  PIN out2[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 144.530 486.220 144.810 490.220 ;
    END
  END out2[20]
  PIN out2[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END out2[21]
  PIN out2[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 477.400 479.500 478.000 ;
    END
  END out2[22]
  PIN out2[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END out2[23]
  PIN out2[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 225.800 479.500 226.400 ;
    END
  END out2[24]
  PIN out2[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END out2[25]
  PIN out2[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 44.920 479.500 45.520 ;
    END
  END out2[26]
  PIN out2[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END out2[27]
  PIN out2[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 427.890 486.220 428.170 490.220 ;
    END
  END out2[28]
  PIN out2[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END out2[29]
  PIN out2[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 232.850 486.220 233.130 490.220 ;
    END
  END out2[2]
  PIN out2[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END out2[30]
  PIN out2[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END out2[31]
  PIN out2[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.730 486.220 62.010 490.220 ;
    END
  END out2[3]
  PIN out2[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.130 486.220 379.410 490.220 ;
    END
  END out2[4]
  PIN out2[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 184.090 486.220 184.370 490.220 ;
    END
  END out2[5]
  PIN out2[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END out2[6]
  PIN out2[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 188.690 486.220 188.970 490.220 ;
    END
  END out2[7]
  PIN out2[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END out2[8]
  PIN out2[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 59.880 479.500 60.480 ;
    END
  END out2[9]
  PIN out3[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END out3[0]
  PIN out3[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 422.370 486.220 422.650 490.220 ;
    END
  END out3[10]
  PIN out3[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 271.490 486.220 271.770 490.220 ;
    END
  END out3[11]
  PIN out3[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 339.570 486.220 339.850 490.220 ;
    END
  END out3[12]
  PIN out3[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END out3[13]
  PIN out3[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END out3[14]
  PIN out3[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 276.120 479.500 276.720 ;
    END
  END out3[15]
  PIN out3[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END out3[16]
  PIN out3[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END out3[17]
  PIN out3[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 349.690 486.220 349.970 490.220 ;
    END
  END out3[18]
  PIN out3[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.170 486.220 91.450 490.220 ;
    END
  END out3[19]
  PIN out3[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 57.130 486.220 57.410 490.220 ;
    END
  END out3[1]
  PIN out3[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END out3[20]
  PIN out3[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END out3[21]
  PIN out3[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END out3[22]
  PIN out3[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 256.770 486.220 257.050 490.220 ;
    END
  END out3[23]
  PIN out3[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END out3[24]
  PIN out3[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 81.640 479.500 82.240 ;
    END
  END out3[25]
  PIN out3[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END out3[26]
  PIN out3[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 486.220 8.650 490.220 ;
    END
  END out3[27]
  PIN out3[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.290 486.220 354.570 490.220 ;
    END
  END out3[28]
  PIN out3[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.930 486.220 393.210 490.220 ;
    END
  END out3[29]
  PIN out3[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END out3[2]
  PIN out3[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END out3[30]
  PIN out3[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END out3[31]
  PIN out3[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END out3[3]
  PIN out3[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END out3[4]
  PIN out3[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.730 486.220 223.010 490.220 ;
    END
  END out3[5]
  PIN out3[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END out3[6]
  PIN out3[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.500 9.560 479.500 10.160 ;
    END
  END out3[7]
  PIN out3[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END out3[8]
  PIN out3[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 471.130 486.220 471.410 490.220 ;
    END
  END out3[9]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END rst
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 473.800 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 473.800 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 473.800 478.805 ;
      LAYER met1 ;
        RECT 2.830 4.460 476.030 483.100 ;
      LAYER met2 ;
        RECT 2.860 485.940 3.490 486.220 ;
        RECT 4.330 485.940 8.090 486.220 ;
        RECT 8.930 485.940 12.690 486.220 ;
        RECT 13.530 485.940 17.290 486.220 ;
        RECT 18.130 485.940 22.810 486.220 ;
        RECT 23.650 485.940 27.410 486.220 ;
        RECT 28.250 485.940 32.010 486.220 ;
        RECT 32.850 485.940 37.530 486.220 ;
        RECT 38.370 485.940 42.130 486.220 ;
        RECT 42.970 485.940 46.730 486.220 ;
        RECT 47.570 485.940 52.250 486.220 ;
        RECT 53.090 485.940 56.850 486.220 ;
        RECT 57.690 485.940 61.450 486.220 ;
        RECT 62.290 485.940 66.050 486.220 ;
        RECT 66.890 485.940 71.570 486.220 ;
        RECT 72.410 485.940 76.170 486.220 ;
        RECT 77.010 485.940 80.770 486.220 ;
        RECT 81.610 485.940 86.290 486.220 ;
        RECT 87.130 485.940 90.890 486.220 ;
        RECT 91.730 485.940 95.490 486.220 ;
        RECT 96.330 485.940 100.090 486.220 ;
        RECT 100.930 485.940 105.610 486.220 ;
        RECT 106.450 485.940 110.210 486.220 ;
        RECT 111.050 485.940 114.810 486.220 ;
        RECT 115.650 485.940 120.330 486.220 ;
        RECT 121.170 485.940 124.930 486.220 ;
        RECT 125.770 485.940 129.530 486.220 ;
        RECT 130.370 485.940 135.050 486.220 ;
        RECT 135.890 485.940 139.650 486.220 ;
        RECT 140.490 485.940 144.250 486.220 ;
        RECT 145.090 485.940 148.850 486.220 ;
        RECT 149.690 485.940 154.370 486.220 ;
        RECT 155.210 485.940 158.970 486.220 ;
        RECT 159.810 485.940 163.570 486.220 ;
        RECT 164.410 485.940 169.090 486.220 ;
        RECT 169.930 485.940 173.690 486.220 ;
        RECT 174.530 485.940 178.290 486.220 ;
        RECT 179.130 485.940 183.810 486.220 ;
        RECT 184.650 485.940 188.410 486.220 ;
        RECT 189.250 485.940 193.010 486.220 ;
        RECT 193.850 485.940 197.610 486.220 ;
        RECT 198.450 485.940 203.130 486.220 ;
        RECT 203.970 485.940 207.730 486.220 ;
        RECT 208.570 485.940 212.330 486.220 ;
        RECT 213.170 485.940 217.850 486.220 ;
        RECT 218.690 485.940 222.450 486.220 ;
        RECT 223.290 485.940 227.050 486.220 ;
        RECT 227.890 485.940 232.570 486.220 ;
        RECT 233.410 485.940 237.170 486.220 ;
        RECT 238.010 485.940 241.770 486.220 ;
        RECT 242.610 485.940 246.370 486.220 ;
        RECT 247.210 485.940 251.890 486.220 ;
        RECT 252.730 485.940 256.490 486.220 ;
        RECT 257.330 485.940 261.090 486.220 ;
        RECT 261.930 485.940 266.610 486.220 ;
        RECT 267.450 485.940 271.210 486.220 ;
        RECT 272.050 485.940 275.810 486.220 ;
        RECT 276.650 485.940 281.330 486.220 ;
        RECT 282.170 485.940 285.930 486.220 ;
        RECT 286.770 485.940 290.530 486.220 ;
        RECT 291.370 485.940 295.130 486.220 ;
        RECT 295.970 485.940 300.650 486.220 ;
        RECT 301.490 485.940 305.250 486.220 ;
        RECT 306.090 485.940 309.850 486.220 ;
        RECT 310.690 485.940 315.370 486.220 ;
        RECT 316.210 485.940 319.970 486.220 ;
        RECT 320.810 485.940 324.570 486.220 ;
        RECT 325.410 485.940 330.090 486.220 ;
        RECT 330.930 485.940 334.690 486.220 ;
        RECT 335.530 485.940 339.290 486.220 ;
        RECT 340.130 485.940 343.890 486.220 ;
        RECT 344.730 485.940 349.410 486.220 ;
        RECT 350.250 485.940 354.010 486.220 ;
        RECT 354.850 485.940 358.610 486.220 ;
        RECT 359.450 485.940 364.130 486.220 ;
        RECT 364.970 485.940 368.730 486.220 ;
        RECT 369.570 485.940 373.330 486.220 ;
        RECT 374.170 485.940 378.850 486.220 ;
        RECT 379.690 485.940 383.450 486.220 ;
        RECT 384.290 485.940 388.050 486.220 ;
        RECT 388.890 485.940 392.650 486.220 ;
        RECT 393.490 485.940 398.170 486.220 ;
        RECT 399.010 485.940 402.770 486.220 ;
        RECT 403.610 485.940 407.370 486.220 ;
        RECT 408.210 485.940 412.890 486.220 ;
        RECT 413.730 485.940 417.490 486.220 ;
        RECT 418.330 485.940 422.090 486.220 ;
        RECT 422.930 485.940 427.610 486.220 ;
        RECT 428.450 485.940 432.210 486.220 ;
        RECT 433.050 485.940 436.810 486.220 ;
        RECT 437.650 485.940 441.410 486.220 ;
        RECT 442.250 485.940 446.930 486.220 ;
        RECT 447.770 485.940 451.530 486.220 ;
        RECT 452.370 485.940 456.130 486.220 ;
        RECT 456.970 485.940 461.650 486.220 ;
        RECT 462.490 485.940 466.250 486.220 ;
        RECT 467.090 485.940 470.850 486.220 ;
        RECT 471.690 485.940 475.450 486.220 ;
        RECT 2.860 4.280 476.000 485.940 ;
        RECT 3.410 4.000 7.170 4.280 ;
        RECT 8.010 4.000 11.770 4.280 ;
        RECT 12.610 4.000 16.370 4.280 ;
        RECT 17.210 4.000 21.890 4.280 ;
        RECT 22.730 4.000 26.490 4.280 ;
        RECT 27.330 4.000 31.090 4.280 ;
        RECT 31.930 4.000 36.610 4.280 ;
        RECT 37.450 4.000 41.210 4.280 ;
        RECT 42.050 4.000 45.810 4.280 ;
        RECT 46.650 4.000 50.410 4.280 ;
        RECT 51.250 4.000 55.930 4.280 ;
        RECT 56.770 4.000 60.530 4.280 ;
        RECT 61.370 4.000 65.130 4.280 ;
        RECT 65.970 4.000 70.650 4.280 ;
        RECT 71.490 4.000 75.250 4.280 ;
        RECT 76.090 4.000 79.850 4.280 ;
        RECT 80.690 4.000 85.370 4.280 ;
        RECT 86.210 4.000 89.970 4.280 ;
        RECT 90.810 4.000 94.570 4.280 ;
        RECT 95.410 4.000 99.170 4.280 ;
        RECT 100.010 4.000 104.690 4.280 ;
        RECT 105.530 4.000 109.290 4.280 ;
        RECT 110.130 4.000 113.890 4.280 ;
        RECT 114.730 4.000 119.410 4.280 ;
        RECT 120.250 4.000 124.010 4.280 ;
        RECT 124.850 4.000 128.610 4.280 ;
        RECT 129.450 4.000 134.130 4.280 ;
        RECT 134.970 4.000 138.730 4.280 ;
        RECT 139.570 4.000 143.330 4.280 ;
        RECT 144.170 4.000 147.930 4.280 ;
        RECT 148.770 4.000 153.450 4.280 ;
        RECT 154.290 4.000 158.050 4.280 ;
        RECT 158.890 4.000 162.650 4.280 ;
        RECT 163.490 4.000 168.170 4.280 ;
        RECT 169.010 4.000 172.770 4.280 ;
        RECT 173.610 4.000 177.370 4.280 ;
        RECT 178.210 4.000 182.890 4.280 ;
        RECT 183.730 4.000 187.490 4.280 ;
        RECT 188.330 4.000 192.090 4.280 ;
        RECT 192.930 4.000 196.690 4.280 ;
        RECT 197.530 4.000 202.210 4.280 ;
        RECT 203.050 4.000 206.810 4.280 ;
        RECT 207.650 4.000 211.410 4.280 ;
        RECT 212.250 4.000 216.930 4.280 ;
        RECT 217.770 4.000 221.530 4.280 ;
        RECT 222.370 4.000 226.130 4.280 ;
        RECT 226.970 4.000 231.650 4.280 ;
        RECT 232.490 4.000 236.250 4.280 ;
        RECT 237.090 4.000 240.850 4.280 ;
        RECT 241.690 4.000 245.450 4.280 ;
        RECT 246.290 4.000 250.970 4.280 ;
        RECT 251.810 4.000 255.570 4.280 ;
        RECT 256.410 4.000 260.170 4.280 ;
        RECT 261.010 4.000 265.690 4.280 ;
        RECT 266.530 4.000 270.290 4.280 ;
        RECT 271.130 4.000 274.890 4.280 ;
        RECT 275.730 4.000 280.410 4.280 ;
        RECT 281.250 4.000 285.010 4.280 ;
        RECT 285.850 4.000 289.610 4.280 ;
        RECT 290.450 4.000 294.210 4.280 ;
        RECT 295.050 4.000 299.730 4.280 ;
        RECT 300.570 4.000 304.330 4.280 ;
        RECT 305.170 4.000 308.930 4.280 ;
        RECT 309.770 4.000 314.450 4.280 ;
        RECT 315.290 4.000 319.050 4.280 ;
        RECT 319.890 4.000 323.650 4.280 ;
        RECT 324.490 4.000 329.170 4.280 ;
        RECT 330.010 4.000 333.770 4.280 ;
        RECT 334.610 4.000 338.370 4.280 ;
        RECT 339.210 4.000 342.970 4.280 ;
        RECT 343.810 4.000 348.490 4.280 ;
        RECT 349.330 4.000 353.090 4.280 ;
        RECT 353.930 4.000 357.690 4.280 ;
        RECT 358.530 4.000 363.210 4.280 ;
        RECT 364.050 4.000 367.810 4.280 ;
        RECT 368.650 4.000 372.410 4.280 ;
        RECT 373.250 4.000 377.930 4.280 ;
        RECT 378.770 4.000 382.530 4.280 ;
        RECT 383.370 4.000 387.130 4.280 ;
        RECT 387.970 4.000 391.730 4.280 ;
        RECT 392.570 4.000 397.250 4.280 ;
        RECT 398.090 4.000 401.850 4.280 ;
        RECT 402.690 4.000 406.450 4.280 ;
        RECT 407.290 4.000 411.970 4.280 ;
        RECT 412.810 4.000 416.570 4.280 ;
        RECT 417.410 4.000 421.170 4.280 ;
        RECT 422.010 4.000 425.770 4.280 ;
        RECT 426.610 4.000 431.290 4.280 ;
        RECT 432.130 4.000 435.890 4.280 ;
        RECT 436.730 4.000 440.490 4.280 ;
        RECT 441.330 4.000 446.010 4.280 ;
        RECT 446.850 4.000 450.610 4.280 ;
        RECT 451.450 4.000 455.210 4.280 ;
        RECT 456.050 4.000 460.730 4.280 ;
        RECT 461.570 4.000 465.330 4.280 ;
        RECT 466.170 4.000 469.930 4.280 ;
        RECT 470.770 4.000 474.530 4.280 ;
        RECT 475.370 4.000 476.000 4.280 ;
      LAYER met3 ;
        RECT 4.000 479.760 475.500 486.025 ;
        RECT 4.400 478.400 475.500 479.760 ;
        RECT 4.400 478.360 475.100 478.400 ;
        RECT 4.000 477.000 475.100 478.360 ;
        RECT 4.000 472.960 475.500 477.000 ;
        RECT 4.400 471.600 475.500 472.960 ;
        RECT 4.400 471.560 475.100 471.600 ;
        RECT 4.000 470.200 475.100 471.560 ;
        RECT 4.000 466.160 475.500 470.200 ;
        RECT 4.400 464.800 475.500 466.160 ;
        RECT 4.400 464.760 475.100 464.800 ;
        RECT 4.000 463.400 475.100 464.760 ;
        RECT 4.000 458.000 475.500 463.400 ;
        RECT 4.400 456.640 475.500 458.000 ;
        RECT 4.400 456.600 475.100 456.640 ;
        RECT 4.000 455.240 475.100 456.600 ;
        RECT 4.000 451.200 475.500 455.240 ;
        RECT 4.400 449.840 475.500 451.200 ;
        RECT 4.400 449.800 475.100 449.840 ;
        RECT 4.000 448.440 475.100 449.800 ;
        RECT 4.000 444.400 475.500 448.440 ;
        RECT 4.400 443.040 475.500 444.400 ;
        RECT 4.400 443.000 475.100 443.040 ;
        RECT 4.000 441.640 475.100 443.000 ;
        RECT 4.000 436.240 475.500 441.640 ;
        RECT 4.400 434.880 475.500 436.240 ;
        RECT 4.400 434.840 475.100 434.880 ;
        RECT 4.000 433.480 475.100 434.840 ;
        RECT 4.000 429.440 475.500 433.480 ;
        RECT 4.400 428.080 475.500 429.440 ;
        RECT 4.400 428.040 475.100 428.080 ;
        RECT 4.000 426.680 475.100 428.040 ;
        RECT 4.000 422.640 475.500 426.680 ;
        RECT 4.400 421.280 475.500 422.640 ;
        RECT 4.400 421.240 475.100 421.280 ;
        RECT 4.000 419.880 475.100 421.240 ;
        RECT 4.000 415.840 475.500 419.880 ;
        RECT 4.400 414.480 475.500 415.840 ;
        RECT 4.400 414.440 475.100 414.480 ;
        RECT 4.000 413.080 475.100 414.440 ;
        RECT 4.000 407.680 475.500 413.080 ;
        RECT 4.400 406.320 475.500 407.680 ;
        RECT 4.400 406.280 475.100 406.320 ;
        RECT 4.000 404.920 475.100 406.280 ;
        RECT 4.000 400.880 475.500 404.920 ;
        RECT 4.400 399.520 475.500 400.880 ;
        RECT 4.400 399.480 475.100 399.520 ;
        RECT 4.000 398.120 475.100 399.480 ;
        RECT 4.000 394.080 475.500 398.120 ;
        RECT 4.400 392.720 475.500 394.080 ;
        RECT 4.400 392.680 475.100 392.720 ;
        RECT 4.000 391.320 475.100 392.680 ;
        RECT 4.000 385.920 475.500 391.320 ;
        RECT 4.400 384.560 475.500 385.920 ;
        RECT 4.400 384.520 475.100 384.560 ;
        RECT 4.000 383.160 475.100 384.520 ;
        RECT 4.000 379.120 475.500 383.160 ;
        RECT 4.400 377.760 475.500 379.120 ;
        RECT 4.400 377.720 475.100 377.760 ;
        RECT 4.000 376.360 475.100 377.720 ;
        RECT 4.000 372.320 475.500 376.360 ;
        RECT 4.400 370.960 475.500 372.320 ;
        RECT 4.400 370.920 475.100 370.960 ;
        RECT 4.000 369.560 475.100 370.920 ;
        RECT 4.000 364.160 475.500 369.560 ;
        RECT 4.400 362.800 475.500 364.160 ;
        RECT 4.400 362.760 475.100 362.800 ;
        RECT 4.000 361.400 475.100 362.760 ;
        RECT 4.000 357.360 475.500 361.400 ;
        RECT 4.400 356.000 475.500 357.360 ;
        RECT 4.400 355.960 475.100 356.000 ;
        RECT 4.000 354.600 475.100 355.960 ;
        RECT 4.000 350.560 475.500 354.600 ;
        RECT 4.400 349.200 475.500 350.560 ;
        RECT 4.400 349.160 475.100 349.200 ;
        RECT 4.000 347.800 475.100 349.160 ;
        RECT 4.000 343.760 475.500 347.800 ;
        RECT 4.400 342.400 475.500 343.760 ;
        RECT 4.400 342.360 475.100 342.400 ;
        RECT 4.000 341.000 475.100 342.360 ;
        RECT 4.000 335.600 475.500 341.000 ;
        RECT 4.400 334.240 475.500 335.600 ;
        RECT 4.400 334.200 475.100 334.240 ;
        RECT 4.000 332.840 475.100 334.200 ;
        RECT 4.000 328.800 475.500 332.840 ;
        RECT 4.400 327.440 475.500 328.800 ;
        RECT 4.400 327.400 475.100 327.440 ;
        RECT 4.000 326.040 475.100 327.400 ;
        RECT 4.000 322.000 475.500 326.040 ;
        RECT 4.400 320.640 475.500 322.000 ;
        RECT 4.400 320.600 475.100 320.640 ;
        RECT 4.000 319.240 475.100 320.600 ;
        RECT 4.000 313.840 475.500 319.240 ;
        RECT 4.400 312.480 475.500 313.840 ;
        RECT 4.400 312.440 475.100 312.480 ;
        RECT 4.000 311.080 475.100 312.440 ;
        RECT 4.000 307.040 475.500 311.080 ;
        RECT 4.400 305.680 475.500 307.040 ;
        RECT 4.400 305.640 475.100 305.680 ;
        RECT 4.000 304.280 475.100 305.640 ;
        RECT 4.000 300.240 475.500 304.280 ;
        RECT 4.400 298.880 475.500 300.240 ;
        RECT 4.400 298.840 475.100 298.880 ;
        RECT 4.000 297.480 475.100 298.840 ;
        RECT 4.000 292.080 475.500 297.480 ;
        RECT 4.400 290.720 475.500 292.080 ;
        RECT 4.400 290.680 475.100 290.720 ;
        RECT 4.000 289.320 475.100 290.680 ;
        RECT 4.000 285.280 475.500 289.320 ;
        RECT 4.400 283.920 475.500 285.280 ;
        RECT 4.400 283.880 475.100 283.920 ;
        RECT 4.000 282.520 475.100 283.880 ;
        RECT 4.000 278.480 475.500 282.520 ;
        RECT 4.400 277.120 475.500 278.480 ;
        RECT 4.400 277.080 475.100 277.120 ;
        RECT 4.000 275.720 475.100 277.080 ;
        RECT 4.000 271.680 475.500 275.720 ;
        RECT 4.400 270.320 475.500 271.680 ;
        RECT 4.400 270.280 475.100 270.320 ;
        RECT 4.000 268.920 475.100 270.280 ;
        RECT 4.000 263.520 475.500 268.920 ;
        RECT 4.400 262.160 475.500 263.520 ;
        RECT 4.400 262.120 475.100 262.160 ;
        RECT 4.000 260.760 475.100 262.120 ;
        RECT 4.000 256.720 475.500 260.760 ;
        RECT 4.400 255.360 475.500 256.720 ;
        RECT 4.400 255.320 475.100 255.360 ;
        RECT 4.000 253.960 475.100 255.320 ;
        RECT 4.000 249.920 475.500 253.960 ;
        RECT 4.400 248.560 475.500 249.920 ;
        RECT 4.400 248.520 475.100 248.560 ;
        RECT 4.000 247.160 475.100 248.520 ;
        RECT 4.000 241.760 475.500 247.160 ;
        RECT 4.400 240.400 475.500 241.760 ;
        RECT 4.400 240.360 475.100 240.400 ;
        RECT 4.000 239.000 475.100 240.360 ;
        RECT 4.000 234.960 475.500 239.000 ;
        RECT 4.400 233.600 475.500 234.960 ;
        RECT 4.400 233.560 475.100 233.600 ;
        RECT 4.000 232.200 475.100 233.560 ;
        RECT 4.000 228.160 475.500 232.200 ;
        RECT 4.400 226.800 475.500 228.160 ;
        RECT 4.400 226.760 475.100 226.800 ;
        RECT 4.000 225.400 475.100 226.760 ;
        RECT 4.000 220.000 475.500 225.400 ;
        RECT 4.400 218.640 475.500 220.000 ;
        RECT 4.400 218.600 475.100 218.640 ;
        RECT 4.000 217.240 475.100 218.600 ;
        RECT 4.000 213.200 475.500 217.240 ;
        RECT 4.400 211.840 475.500 213.200 ;
        RECT 4.400 211.800 475.100 211.840 ;
        RECT 4.000 210.440 475.100 211.800 ;
        RECT 4.000 206.400 475.500 210.440 ;
        RECT 4.400 205.040 475.500 206.400 ;
        RECT 4.400 205.000 475.100 205.040 ;
        RECT 4.000 203.640 475.100 205.000 ;
        RECT 4.000 199.600 475.500 203.640 ;
        RECT 4.400 198.240 475.500 199.600 ;
        RECT 4.400 198.200 475.100 198.240 ;
        RECT 4.000 196.840 475.100 198.200 ;
        RECT 4.000 191.440 475.500 196.840 ;
        RECT 4.400 190.080 475.500 191.440 ;
        RECT 4.400 190.040 475.100 190.080 ;
        RECT 4.000 188.680 475.100 190.040 ;
        RECT 4.000 184.640 475.500 188.680 ;
        RECT 4.400 183.280 475.500 184.640 ;
        RECT 4.400 183.240 475.100 183.280 ;
        RECT 4.000 181.880 475.100 183.240 ;
        RECT 4.000 177.840 475.500 181.880 ;
        RECT 4.400 176.480 475.500 177.840 ;
        RECT 4.400 176.440 475.100 176.480 ;
        RECT 4.000 175.080 475.100 176.440 ;
        RECT 4.000 169.680 475.500 175.080 ;
        RECT 4.400 168.320 475.500 169.680 ;
        RECT 4.400 168.280 475.100 168.320 ;
        RECT 4.000 166.920 475.100 168.280 ;
        RECT 4.000 162.880 475.500 166.920 ;
        RECT 4.400 161.520 475.500 162.880 ;
        RECT 4.400 161.480 475.100 161.520 ;
        RECT 4.000 160.120 475.100 161.480 ;
        RECT 4.000 156.080 475.500 160.120 ;
        RECT 4.400 154.720 475.500 156.080 ;
        RECT 4.400 154.680 475.100 154.720 ;
        RECT 4.000 153.320 475.100 154.680 ;
        RECT 4.000 147.920 475.500 153.320 ;
        RECT 4.400 146.560 475.500 147.920 ;
        RECT 4.400 146.520 475.100 146.560 ;
        RECT 4.000 145.160 475.100 146.520 ;
        RECT 4.000 141.120 475.500 145.160 ;
        RECT 4.400 139.760 475.500 141.120 ;
        RECT 4.400 139.720 475.100 139.760 ;
        RECT 4.000 138.360 475.100 139.720 ;
        RECT 4.000 134.320 475.500 138.360 ;
        RECT 4.400 132.960 475.500 134.320 ;
        RECT 4.400 132.920 475.100 132.960 ;
        RECT 4.000 131.560 475.100 132.920 ;
        RECT 4.000 127.520 475.500 131.560 ;
        RECT 4.400 126.160 475.500 127.520 ;
        RECT 4.400 126.120 475.100 126.160 ;
        RECT 4.000 124.760 475.100 126.120 ;
        RECT 4.000 119.360 475.500 124.760 ;
        RECT 4.400 118.000 475.500 119.360 ;
        RECT 4.400 117.960 475.100 118.000 ;
        RECT 4.000 116.600 475.100 117.960 ;
        RECT 4.000 112.560 475.500 116.600 ;
        RECT 4.400 111.200 475.500 112.560 ;
        RECT 4.400 111.160 475.100 111.200 ;
        RECT 4.000 109.800 475.100 111.160 ;
        RECT 4.000 105.760 475.500 109.800 ;
        RECT 4.400 104.400 475.500 105.760 ;
        RECT 4.400 104.360 475.100 104.400 ;
        RECT 4.000 103.000 475.100 104.360 ;
        RECT 4.000 97.600 475.500 103.000 ;
        RECT 4.400 96.240 475.500 97.600 ;
        RECT 4.400 96.200 475.100 96.240 ;
        RECT 4.000 94.840 475.100 96.200 ;
        RECT 4.000 90.800 475.500 94.840 ;
        RECT 4.400 89.440 475.500 90.800 ;
        RECT 4.400 89.400 475.100 89.440 ;
        RECT 4.000 88.040 475.100 89.400 ;
        RECT 4.000 84.000 475.500 88.040 ;
        RECT 4.400 82.640 475.500 84.000 ;
        RECT 4.400 82.600 475.100 82.640 ;
        RECT 4.000 81.240 475.100 82.600 ;
        RECT 4.000 75.840 475.500 81.240 ;
        RECT 4.400 74.480 475.500 75.840 ;
        RECT 4.400 74.440 475.100 74.480 ;
        RECT 4.000 73.080 475.100 74.440 ;
        RECT 4.000 69.040 475.500 73.080 ;
        RECT 4.400 67.680 475.500 69.040 ;
        RECT 4.400 67.640 475.100 67.680 ;
        RECT 4.000 66.280 475.100 67.640 ;
        RECT 4.000 62.240 475.500 66.280 ;
        RECT 4.400 60.880 475.500 62.240 ;
        RECT 4.400 60.840 475.100 60.880 ;
        RECT 4.000 59.480 475.100 60.840 ;
        RECT 4.000 55.440 475.500 59.480 ;
        RECT 4.400 54.080 475.500 55.440 ;
        RECT 4.400 54.040 475.100 54.080 ;
        RECT 4.000 52.680 475.100 54.040 ;
        RECT 4.000 47.280 475.500 52.680 ;
        RECT 4.400 45.920 475.500 47.280 ;
        RECT 4.400 45.880 475.100 45.920 ;
        RECT 4.000 44.520 475.100 45.880 ;
        RECT 4.000 40.480 475.500 44.520 ;
        RECT 4.400 39.120 475.500 40.480 ;
        RECT 4.400 39.080 475.100 39.120 ;
        RECT 4.000 37.720 475.100 39.080 ;
        RECT 4.000 33.680 475.500 37.720 ;
        RECT 4.400 32.320 475.500 33.680 ;
        RECT 4.400 32.280 475.100 32.320 ;
        RECT 4.000 30.920 475.100 32.280 ;
        RECT 4.000 25.520 475.500 30.920 ;
        RECT 4.400 24.160 475.500 25.520 ;
        RECT 4.400 24.120 475.100 24.160 ;
        RECT 4.000 22.760 475.100 24.120 ;
        RECT 4.000 18.720 475.500 22.760 ;
        RECT 4.400 17.360 475.500 18.720 ;
        RECT 4.400 17.320 475.100 17.360 ;
        RECT 4.000 15.960 475.100 17.320 ;
        RECT 4.000 11.920 475.500 15.960 ;
        RECT 4.400 10.560 475.500 11.920 ;
        RECT 4.400 10.520 475.100 10.560 ;
        RECT 4.000 9.695 475.100 10.520 ;
      LAYER met4 ;
        RECT 16.855 10.640 458.785 478.960 ;
      LAYER met5 ;
        RECT 5.520 179.670 473.800 411.040 ;
  END
END mac_cluster
END LIBRARY

