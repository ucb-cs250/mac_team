VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mac_cluster
  CLASS BLOCK ;
  FOREIGN mac_cluster ;
  ORIGIN 0.000 0.000 ;
  SIZE 499.950 BY 510.670 ;
  PIN A0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.850 506.670 187.130 510.670 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 273.400 499.950 274.000 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 4.000 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 420.530 506.670 420.810 510.670 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 201.570 506.670 201.850 510.670 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END A0[7]
  PIN A1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.730 506.670 177.010 510.670 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 469.240 499.950 469.840 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.210 506.670 263.490 510.670 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.050 506.670 288.330 510.670 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 506.670 18.770 510.670 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 273.330 506.670 273.610 510.670 ;
    END
  END A1[7]
  PIN A2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 451.810 506.670 452.090 510.670 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END A2[6]
  PIN A2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 446.120 499.950 446.720 ;
    END
  END A2[7]
  PIN A3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 237.450 506.670 237.730 510.670 ;
    END
  END A3[0]
  PIN A3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END A3[1]
  PIN A3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 466.530 506.670 466.810 510.670 ;
    END
  END A3[2]
  PIN A3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 207.090 506.670 207.370 510.670 ;
    END
  END A3[3]
  PIN A3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END A3[4]
  PIN A3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END A3[5]
  PIN A3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END A3[6]
  PIN A3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.090 506.670 69.370 510.670 ;
    END
  END A3[7]
  PIN B0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END B0[0]
  PIN B0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END B0[1]
  PIN B0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END B0[2]
  PIN B0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END B0[3]
  PIN B0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 220.360 499.950 220.960 ;
    END
  END B0[4]
  PIN B0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.330 506.670 227.610 510.670 ;
    END
  END B0[5]
  PIN B0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 506.670 74.890 510.670 ;
    END
  END B0[6]
  PIN B0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END B0[7]
  PIN B1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.450 506.670 145.730 510.670 ;
    END
  END B1[0]
  PIN B1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 371.320 499.950 371.920 ;
    END
  END B1[1]
  PIN B1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 152.360 499.950 152.960 ;
    END
  END B1[2]
  PIN B1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END B1[3]
  PIN B1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 375.450 506.670 375.730 510.670 ;
    END
  END B1[4]
  PIN B1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END B1[5]
  PIN B1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.490 506.670 156.770 510.670 ;
    END
  END B1[6]
  PIN B1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 243.480 499.950 244.080 ;
    END
  END B1[7]
  PIN B2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END B2[0]
  PIN B2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END B2[1]
  PIN B2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END B2[2]
  PIN B2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 115.640 499.950 116.240 ;
    END
  END B2[3]
  PIN B2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 161.090 506.670 161.370 510.670 ;
    END
  END B2[4]
  PIN B2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 506.670 24.290 510.670 ;
    END
  END B2[5]
  PIN B2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END B2[6]
  PIN B2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 280.200 499.950 280.800 ;
    END
  END B2[7]
  PIN B3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 77.560 499.950 78.160 ;
    END
  END B3[0]
  PIN B3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END B3[1]
  PIN B3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END B3[2]
  PIN B3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 484.200 499.950 484.800 ;
    END
  END B3[3]
  PIN B3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 213.560 499.950 214.160 ;
    END
  END B3[4]
  PIN B3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 506.670 28.890 510.670 ;
    END
  END B3[5]
  PIN B3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END B3[6]
  PIN B3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 107.480 499.950 108.080 ;
    END
  END B3[7]
  PIN cfg[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 257.690 506.670 257.970 510.670 ;
    END
  END cfg[0]
  PIN cfg[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END cfg[100]
  PIN cfg[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END cfg[101]
  PIN cfg[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END cfg[102]
  PIN cfg[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 506.670 49.130 510.670 ;
    END
  END cfg[103]
  PIN cfg[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END cfg[104]
  PIN cfg[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END cfg[105]
  PIN cfg[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 431.160 499.950 431.760 ;
    END
  END cfg[106]
  PIN cfg[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END cfg[107]
  PIN cfg[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END cfg[108]
  PIN cfg[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 506.670 110.770 510.670 ;
    END
  END cfg[109]
  PIN cfg[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END cfg[10]
  PIN cfg[110]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END cfg[110]
  PIN cfg[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END cfg[111]
  PIN cfg[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END cfg[112]
  PIN cfg[113]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 205.400 499.950 206.000 ;
    END
  END cfg[113]
  PIN cfg[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 250.280 499.950 250.880 ;
    END
  END cfg[114]
  PIN cfg[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.250 506.670 90.530 510.670 ;
    END
  END cfg[115]
  PIN cfg[116]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END cfg[116]
  PIN cfg[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 431.570 506.670 431.850 510.670 ;
    END
  END cfg[117]
  PIN cfg[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END cfg[118]
  PIN cfg[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END cfg[119]
  PIN cfg[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END cfg[11]
  PIN cfg[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 120.610 506.670 120.890 510.670 ;
    END
  END cfg[120]
  PIN cfg[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 24.520 499.950 25.120 ;
    END
  END cfg[121]
  PIN cfg[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END cfg[122]
  PIN cfg[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END cfg[123]
  PIN cfg[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 363.160 499.950 363.760 ;
    END
  END cfg[124]
  PIN cfg[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 506.670 34.410 510.670 ;
    END
  END cfg[125]
  PIN cfg[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 258.440 499.950 259.040 ;
    END
  END cfg[126]
  PIN cfg[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END cfg[127]
  PIN cfg[128]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END cfg[128]
  PIN cfg[129]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END cfg[129]
  PIN cfg[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END cfg[12]
  PIN cfg[130]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END cfg[130]
  PIN cfg[131]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 349.690 506.670 349.970 510.670 ;
    END
  END cfg[131]
  PIN cfg[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.930 506.670 324.210 510.670 ;
    END
  END cfg[13]
  PIN cfg[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END cfg[14]
  PIN cfg[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END cfg[15]
  PIN cfg[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END cfg[16]
  PIN cfg[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.570 506.670 293.850 510.670 ;
    END
  END cfg[17]
  PIN cfg[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 356.360 499.950 356.960 ;
    END
  END cfg[18]
  PIN cfg[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END cfg[19]
  PIN cfg[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END cfg[1]
  PIN cfg[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 211.690 506.670 211.970 510.670 ;
    END
  END cfg[20]
  PIN cfg[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 92.520 499.950 93.120 ;
    END
  END cfg[21]
  PIN cfg[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 175.480 499.950 176.080 ;
    END
  END cfg[22]
  PIN cfg[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END cfg[23]
  PIN cfg[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 17.720 499.950 18.320 ;
    END
  END cfg[24]
  PIN cfg[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END cfg[25]
  PIN cfg[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END cfg[26]
  PIN cfg[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 339.570 506.670 339.850 510.670 ;
    END
  END cfg[27]
  PIN cfg[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.170 506.670 436.450 510.670 ;
    END
  END cfg[28]
  PIN cfg[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END cfg[29]
  PIN cfg[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END cfg[2]
  PIN cfg[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END cfg[30]
  PIN cfg[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 318.280 499.950 318.880 ;
    END
  END cfg[31]
  PIN cfg[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.050 506.670 472.330 510.670 ;
    END
  END cfg[32]
  PIN cfg[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 253.090 506.670 253.370 510.670 ;
    END
  END cfg[33]
  PIN cfg[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END cfg[34]
  PIN cfg[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END cfg[35]
  PIN cfg[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END cfg[36]
  PIN cfg[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END cfg[37]
  PIN cfg[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 54.440 499.950 55.040 ;
    END
  END cfg[38]
  PIN cfg[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 386.280 499.950 386.880 ;
    END
  END cfg[39]
  PIN cfg[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 461.080 499.950 461.680 ;
    END
  END cfg[3]
  PIN cfg[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END cfg[40]
  PIN cfg[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.730 506.670 85.010 510.670 ;
    END
  END cfg[41]
  PIN cfg[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END cfg[42]
  PIN cfg[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END cfg[43]
  PIN cfg[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 130.600 499.950 131.200 ;
    END
  END cfg[44]
  PIN cfg[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END cfg[45]
  PIN cfg[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 409.400 499.950 410.000 ;
    END
  END cfg[46]
  PIN cfg[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 400.290 506.670 400.570 510.670 ;
    END
  END cfg[47]
  PIN cfg[48]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END cfg[48]
  PIN cfg[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 506.670 79.490 510.670 ;
    END
  END cfg[49]
  PIN cfg[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 171.210 506.670 171.490 510.670 ;
    END
  END cfg[4]
  PIN cfg[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END cfg[50]
  PIN cfg[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.930 506.670 462.210 510.670 ;
    END
  END cfg[51]
  PIN cfg[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END cfg[52]
  PIN cfg[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END cfg[53]
  PIN cfg[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END cfg[54]
  PIN cfg[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END cfg[55]
  PIN cfg[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END cfg[56]
  PIN cfg[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END cfg[57]
  PIN cfg[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 385.570 506.670 385.850 510.670 ;
    END
  END cfg[58]
  PIN cfg[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END cfg[59]
  PIN cfg[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.170 506.670 390.450 510.670 ;
    END
  END cfg[5]
  PIN cfg[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 491.000 499.950 491.600 ;
    END
  END cfg[60]
  PIN cfg[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 295.160 499.950 295.760 ;
    END
  END cfg[61]
  PIN cfg[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.090 506.670 299.370 510.670 ;
    END
  END cfg[62]
  PIN cfg[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 145.560 499.950 146.160 ;
    END
  END cfg[63]
  PIN cfg[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END cfg[64]
  PIN cfg[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END cfg[65]
  PIN cfg[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 506.670 105.250 510.670 ;
    END
  END cfg[66]
  PIN cfg[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 506.670 3.130 510.670 ;
    END
  END cfg[67]
  PIN cfg[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END cfg[68]
  PIN cfg[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END cfg[69]
  PIN cfg[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 303.690 506.670 303.970 510.670 ;
    END
  END cfg[6]
  PIN cfg[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END cfg[70]
  PIN cfg[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 160.520 499.950 161.120 ;
    END
  END cfg[71]
  PIN cfg[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END cfg[72]
  PIN cfg[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END cfg[73]
  PIN cfg[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.610 506.670 166.890 510.670 ;
    END
  END cfg[74]
  PIN cfg[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END cfg[75]
  PIN cfg[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END cfg[76]
  PIN cfg[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END cfg[77]
  PIN cfg[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 32.680 499.950 33.280 ;
    END
  END cfg[78]
  PIN cfg[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 405.810 506.670 406.090 510.670 ;
    END
  END cfg[79]
  PIN cfg[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END cfg[7]
  PIN cfg[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END cfg[80]
  PIN cfg[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END cfg[81]
  PIN cfg[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END cfg[82]
  PIN cfg[83]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END cfg[83]
  PIN cfg[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 505.960 499.950 506.560 ;
    END
  END cfg[84]
  PIN cfg[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 359.810 506.670 360.090 510.670 ;
    END
  END cfg[85]
  PIN cfg[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.330 506.670 319.610 510.670 ;
    END
  END cfg[86]
  PIN cfg[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 198.600 499.950 199.200 ;
    END
  END cfg[87]
  PIN cfg[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.050 506.670 334.330 510.670 ;
    END
  END cfg[88]
  PIN cfg[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END cfg[89]
  PIN cfg[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 333.240 499.950 333.840 ;
    END
  END cfg[8]
  PIN cfg[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END cfg[90]
  PIN cfg[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END cfg[91]
  PIN cfg[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END cfg[92]
  PIN cfg[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END cfg[93]
  PIN cfg[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END cfg[94]
  PIN cfg[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 506.670 115.370 510.670 ;
    END
  END cfg[95]
  PIN cfg[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 100.680 499.950 101.280 ;
    END
  END cfg[96]
  PIN cfg[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END cfg[97]
  PIN cfg[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END cfg[98]
  PIN cfg[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END cfg[99]
  PIN cfg[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 416.200 499.950 416.800 ;
    END
  END cfg[9]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 476.650 506.670 476.930 510.670 ;
    END
  END clk
  PIN cset
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 495.950 228.520 499.950 229.120 ;
    END
  END cset
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 277.930 506.670 278.210 510.670 ;
    END
  END en
  PIN out0[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END out0[0]
  PIN out0[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 415.930 506.670 416.210 510.670 ;
    END
  END out0[10]
  PIN out0[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 265.240 499.950 265.840 ;
    END
  END out0[11]
  PIN out0[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 424.360 499.950 424.960 ;
    END
  END out0[12]
  PIN out0[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 303.320 499.950 303.920 ;
    END
  END out0[13]
  PIN out0[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 122.440 499.950 123.040 ;
    END
  END out0[14]
  PIN out0[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.330 506.670 181.610 510.670 ;
    END
  END out0[15]
  PIN out0[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 140.850 506.670 141.130 510.670 ;
    END
  END out0[16]
  PIN out0[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 125.210 506.670 125.490 510.670 ;
    END
  END out0[17]
  PIN out0[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END out0[18]
  PIN out0[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 415.010 0.000 415.290 4.000 ;
    END
  END out0[19]
  PIN out0[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 341.400 499.950 342.000 ;
    END
  END out0[1]
  PIN out0[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END out0[20]
  PIN out0[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END out0[21]
  PIN out0[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END out0[22]
  PIN out0[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END out0[23]
  PIN out0[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.730 506.670 223.010 510.670 ;
    END
  END out0[24]
  PIN out0[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 380.050 506.670 380.330 510.670 ;
    END
  END out0[25]
  PIN out0[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 401.240 499.950 401.840 ;
    END
  END out0[26]
  PIN out0[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 454.280 499.950 454.880 ;
    END
  END out0[27]
  PIN out0[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.370 506.670 54.650 510.670 ;
    END
  END out0[28]
  PIN out0[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 326.440 499.950 327.040 ;
    END
  END out0[29]
  PIN out0[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 456.410 506.670 456.690 510.670 ;
    END
  END out0[2]
  PIN out0[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END out0[30]
  PIN out0[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END out0[31]
  PIN out0[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END out0[3]
  PIN out0[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 39.480 499.950 40.080 ;
    END
  END out0[4]
  PIN out0[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 378.120 499.950 378.720 ;
    END
  END out0[5]
  PIN out0[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 344.170 506.670 344.450 510.670 ;
    END
  END out0[6]
  PIN out0[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 311.480 499.950 312.080 ;
    END
  END out0[7]
  PIN out0[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END out0[8]
  PIN out0[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 486.770 506.670 487.050 510.670 ;
    END
  END out0[9]
  PIN out1[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 329.450 506.670 329.730 510.670 ;
    END
  END out1[0]
  PIN out1[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 348.200 499.950 348.800 ;
    END
  END out1[10]
  PIN out1[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 439.320 499.950 439.920 ;
    END
  END out1[11]
  PIN out1[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END out1[12]
  PIN out1[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END out1[13]
  PIN out1[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.250 506.670 44.530 510.670 ;
    END
  END out1[14]
  PIN out1[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 309.210 506.670 309.490 510.670 ;
    END
  END out1[15]
  PIN out1[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END out1[16]
  PIN out1[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 190.440 499.950 191.040 ;
    END
  END out1[17]
  PIN out1[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.730 506.670 39.010 510.670 ;
    END
  END out1[18]
  PIN out1[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END out1[19]
  PIN out1[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END out1[1]
  PIN out1[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 476.040 499.950 476.640 ;
    END
  END out1[20]
  PIN out1[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 426.050 506.670 426.330 510.670 ;
    END
  END out1[21]
  PIN out1[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END out1[22]
  PIN out1[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END out1[23]
  PIN out1[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 506.670 131.010 510.670 ;
    END
  END out1[24]
  PIN out1[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END out1[25]
  PIN out1[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END out1[26]
  PIN out1[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 482.170 506.670 482.450 510.670 ;
    END
  END out1[27]
  PIN out1[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 167.320 499.950 167.920 ;
    END
  END out1[28]
  PIN out1[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END out1[29]
  PIN out1[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END out1[2]
  PIN out1[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END out1[30]
  PIN out1[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 506.670 14.170 510.670 ;
    END
  END out1[31]
  PIN out1[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 69.400 499.950 70.000 ;
    END
  END out1[3]
  PIN out1[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END out1[4]
  PIN out1[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END out1[5]
  PIN out1[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END out1[6]
  PIN out1[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 182.280 499.950 182.880 ;
    END
  END out1[7]
  PIN out1[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 217.210 506.670 217.490 510.670 ;
    END
  END out1[8]
  PIN out1[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 506.670 135.610 510.670 ;
    END
  END out1[9]
  PIN out2[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END out2[0]
  PIN out2[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END out2[10]
  PIN out2[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 506.670 100.650 510.670 ;
    END
  END out2[11]
  PIN out2[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 137.400 499.950 138.000 ;
    END
  END out2[12]
  PIN out2[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END out2[13]
  PIN out2[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END out2[14]
  PIN out2[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 247.570 506.670 247.850 510.670 ;
    END
  END out2[15]
  PIN out2[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 313.810 506.670 314.090 510.670 ;
    END
  END out2[16]
  PIN out2[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END out2[17]
  PIN out2[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 393.080 499.950 393.680 ;
    END
  END out2[18]
  PIN out2[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END out2[19]
  PIN out2[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END out2[1]
  PIN out2[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.970 506.670 151.250 510.670 ;
    END
  END out2[20]
  PIN out2[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END out2[21]
  PIN out2[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 499.160 499.950 499.760 ;
    END
  END out2[22]
  PIN out2[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END out2[23]
  PIN out2[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 235.320 499.950 235.920 ;
    END
  END out2[24]
  PIN out2[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END out2[25]
  PIN out2[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 47.640 499.950 48.240 ;
    END
  END out2[26]
  PIN out2[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END out2[27]
  PIN out2[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 446.290 506.670 446.570 510.670 ;
    END
  END out2[28]
  PIN out2[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END out2[29]
  PIN out2[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 242.970 506.670 243.250 510.670 ;
    END
  END out2[2]
  PIN out2[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END out2[30]
  PIN out2[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END out2[31]
  PIN out2[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.490 506.670 64.770 510.670 ;
    END
  END out2[3]
  PIN out2[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.690 506.670 395.970 510.670 ;
    END
  END out2[4]
  PIN out2[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 191.450 506.670 191.730 510.670 ;
    END
  END out2[5]
  PIN out2[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END out2[6]
  PIN out2[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.970 506.670 197.250 510.670 ;
    END
  END out2[7]
  PIN out2[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END out2[8]
  PIN out2[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 62.600 499.950 63.200 ;
    END
  END out2[9]
  PIN out3[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END out3[0]
  PIN out3[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 441.690 506.670 441.970 510.670 ;
    END
  END out3[10]
  PIN out3[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 283.450 506.670 283.730 510.670 ;
    END
  END out3[11]
  PIN out3[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.290 506.670 354.570 510.670 ;
    END
  END out3[12]
  PIN out3[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END out3[13]
  PIN out3[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END out3[14]
  PIN out3[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 288.360 499.950 288.960 ;
    END
  END out3[15]
  PIN out3[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END out3[16]
  PIN out3[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END out3[17]
  PIN out3[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 365.330 506.670 365.610 510.670 ;
    END
  END out3[18]
  PIN out3[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.850 506.670 95.130 510.670 ;
    END
  END out3[19]
  PIN out3[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.970 506.670 59.250 510.670 ;
    END
  END out3[1]
  PIN out3[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END out3[20]
  PIN out3[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END out3[21]
  PIN out3[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END out3[22]
  PIN out3[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 267.810 506.670 268.090 510.670 ;
    END
  END out3[23]
  PIN out3[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END out3[24]
  PIN out3[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 84.360 499.950 84.960 ;
    END
  END out3[25]
  PIN out3[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END out3[26]
  PIN out3[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 506.670 8.650 510.670 ;
    END
  END out3[27]
  PIN out3[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 369.930 506.670 370.210 510.670 ;
    END
  END out3[28]
  PIN out3[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 410.410 506.670 410.690 510.670 ;
    END
  END out3[29]
  PIN out3[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END out3[2]
  PIN out3[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END out3[30]
  PIN out3[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END out3[31]
  PIN out3[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END out3[3]
  PIN out3[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END out3[4]
  PIN out3[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 232.850 506.670 233.130 510.670 ;
    END
  END out3[5]
  PIN out3[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END out3[6]
  PIN out3[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 495.950 9.560 499.950 10.160 ;
    END
  END out3[7]
  PIN out3[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END out3[8]
  PIN out3[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 492.290 506.670 492.570 510.670 ;
    END
  END out3[9]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END rst
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 494.040 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 494.040 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 497.845 ;
      LAYER met1 ;
        RECT 0.070 4.800 497.190 498.740 ;
      LAYER met2 ;
        RECT 0.100 506.390 2.570 506.670 ;
        RECT 3.410 506.390 8.090 506.670 ;
        RECT 8.930 506.390 13.610 506.670 ;
        RECT 14.450 506.390 18.210 506.670 ;
        RECT 19.050 506.390 23.730 506.670 ;
        RECT 24.570 506.390 28.330 506.670 ;
        RECT 29.170 506.390 33.850 506.670 ;
        RECT 34.690 506.390 38.450 506.670 ;
        RECT 39.290 506.390 43.970 506.670 ;
        RECT 44.810 506.390 48.570 506.670 ;
        RECT 49.410 506.390 54.090 506.670 ;
        RECT 54.930 506.390 58.690 506.670 ;
        RECT 59.530 506.390 64.210 506.670 ;
        RECT 65.050 506.390 68.810 506.670 ;
        RECT 69.650 506.390 74.330 506.670 ;
        RECT 75.170 506.390 78.930 506.670 ;
        RECT 79.770 506.390 84.450 506.670 ;
        RECT 85.290 506.390 89.970 506.670 ;
        RECT 90.810 506.390 94.570 506.670 ;
        RECT 95.410 506.390 100.090 506.670 ;
        RECT 100.930 506.390 104.690 506.670 ;
        RECT 105.530 506.390 110.210 506.670 ;
        RECT 111.050 506.390 114.810 506.670 ;
        RECT 115.650 506.390 120.330 506.670 ;
        RECT 121.170 506.390 124.930 506.670 ;
        RECT 125.770 506.390 130.450 506.670 ;
        RECT 131.290 506.390 135.050 506.670 ;
        RECT 135.890 506.390 140.570 506.670 ;
        RECT 141.410 506.390 145.170 506.670 ;
        RECT 146.010 506.390 150.690 506.670 ;
        RECT 151.530 506.390 156.210 506.670 ;
        RECT 157.050 506.390 160.810 506.670 ;
        RECT 161.650 506.390 166.330 506.670 ;
        RECT 167.170 506.390 170.930 506.670 ;
        RECT 171.770 506.390 176.450 506.670 ;
        RECT 177.290 506.390 181.050 506.670 ;
        RECT 181.890 506.390 186.570 506.670 ;
        RECT 187.410 506.390 191.170 506.670 ;
        RECT 192.010 506.390 196.690 506.670 ;
        RECT 197.530 506.390 201.290 506.670 ;
        RECT 202.130 506.390 206.810 506.670 ;
        RECT 207.650 506.390 211.410 506.670 ;
        RECT 212.250 506.390 216.930 506.670 ;
        RECT 217.770 506.390 222.450 506.670 ;
        RECT 223.290 506.390 227.050 506.670 ;
        RECT 227.890 506.390 232.570 506.670 ;
        RECT 233.410 506.390 237.170 506.670 ;
        RECT 238.010 506.390 242.690 506.670 ;
        RECT 243.530 506.390 247.290 506.670 ;
        RECT 248.130 506.390 252.810 506.670 ;
        RECT 253.650 506.390 257.410 506.670 ;
        RECT 258.250 506.390 262.930 506.670 ;
        RECT 263.770 506.390 267.530 506.670 ;
        RECT 268.370 506.390 273.050 506.670 ;
        RECT 273.890 506.390 277.650 506.670 ;
        RECT 278.490 506.390 283.170 506.670 ;
        RECT 284.010 506.390 287.770 506.670 ;
        RECT 288.610 506.390 293.290 506.670 ;
        RECT 294.130 506.390 298.810 506.670 ;
        RECT 299.650 506.390 303.410 506.670 ;
        RECT 304.250 506.390 308.930 506.670 ;
        RECT 309.770 506.390 313.530 506.670 ;
        RECT 314.370 506.390 319.050 506.670 ;
        RECT 319.890 506.390 323.650 506.670 ;
        RECT 324.490 506.390 329.170 506.670 ;
        RECT 330.010 506.390 333.770 506.670 ;
        RECT 334.610 506.390 339.290 506.670 ;
        RECT 340.130 506.390 343.890 506.670 ;
        RECT 344.730 506.390 349.410 506.670 ;
        RECT 350.250 506.390 354.010 506.670 ;
        RECT 354.850 506.390 359.530 506.670 ;
        RECT 360.370 506.390 365.050 506.670 ;
        RECT 365.890 506.390 369.650 506.670 ;
        RECT 370.490 506.390 375.170 506.670 ;
        RECT 376.010 506.390 379.770 506.670 ;
        RECT 380.610 506.390 385.290 506.670 ;
        RECT 386.130 506.390 389.890 506.670 ;
        RECT 390.730 506.390 395.410 506.670 ;
        RECT 396.250 506.390 400.010 506.670 ;
        RECT 400.850 506.390 405.530 506.670 ;
        RECT 406.370 506.390 410.130 506.670 ;
        RECT 410.970 506.390 415.650 506.670 ;
        RECT 416.490 506.390 420.250 506.670 ;
        RECT 421.090 506.390 425.770 506.670 ;
        RECT 426.610 506.390 431.290 506.670 ;
        RECT 432.130 506.390 435.890 506.670 ;
        RECT 436.730 506.390 441.410 506.670 ;
        RECT 442.250 506.390 446.010 506.670 ;
        RECT 446.850 506.390 451.530 506.670 ;
        RECT 452.370 506.390 456.130 506.670 ;
        RECT 456.970 506.390 461.650 506.670 ;
        RECT 462.490 506.390 466.250 506.670 ;
        RECT 467.090 506.390 471.770 506.670 ;
        RECT 472.610 506.390 476.370 506.670 ;
        RECT 477.210 506.390 481.890 506.670 ;
        RECT 482.730 506.390 486.490 506.670 ;
        RECT 487.330 506.390 492.010 506.670 ;
        RECT 492.850 506.390 497.160 506.670 ;
        RECT 0.100 4.280 497.160 506.390 ;
        RECT 0.100 4.000 2.570 4.280 ;
        RECT 3.410 4.000 7.170 4.280 ;
        RECT 8.010 4.000 12.690 4.280 ;
        RECT 13.530 4.000 17.290 4.280 ;
        RECT 18.130 4.000 22.810 4.280 ;
        RECT 23.650 4.000 27.410 4.280 ;
        RECT 28.250 4.000 32.930 4.280 ;
        RECT 33.770 4.000 37.530 4.280 ;
        RECT 38.370 4.000 43.050 4.280 ;
        RECT 43.890 4.000 47.650 4.280 ;
        RECT 48.490 4.000 53.170 4.280 ;
        RECT 54.010 4.000 57.770 4.280 ;
        RECT 58.610 4.000 63.290 4.280 ;
        RECT 64.130 4.000 67.890 4.280 ;
        RECT 68.730 4.000 73.410 4.280 ;
        RECT 74.250 4.000 78.930 4.280 ;
        RECT 79.770 4.000 83.530 4.280 ;
        RECT 84.370 4.000 89.050 4.280 ;
        RECT 89.890 4.000 93.650 4.280 ;
        RECT 94.490 4.000 99.170 4.280 ;
        RECT 100.010 4.000 103.770 4.280 ;
        RECT 104.610 4.000 109.290 4.280 ;
        RECT 110.130 4.000 113.890 4.280 ;
        RECT 114.730 4.000 119.410 4.280 ;
        RECT 120.250 4.000 124.010 4.280 ;
        RECT 124.850 4.000 129.530 4.280 ;
        RECT 130.370 4.000 134.130 4.280 ;
        RECT 134.970 4.000 139.650 4.280 ;
        RECT 140.490 4.000 145.170 4.280 ;
        RECT 146.010 4.000 149.770 4.280 ;
        RECT 150.610 4.000 155.290 4.280 ;
        RECT 156.130 4.000 159.890 4.280 ;
        RECT 160.730 4.000 165.410 4.280 ;
        RECT 166.250 4.000 170.010 4.280 ;
        RECT 170.850 4.000 175.530 4.280 ;
        RECT 176.370 4.000 180.130 4.280 ;
        RECT 180.970 4.000 185.650 4.280 ;
        RECT 186.490 4.000 190.250 4.280 ;
        RECT 191.090 4.000 195.770 4.280 ;
        RECT 196.610 4.000 200.370 4.280 ;
        RECT 201.210 4.000 205.890 4.280 ;
        RECT 206.730 4.000 210.490 4.280 ;
        RECT 211.330 4.000 216.010 4.280 ;
        RECT 216.850 4.000 221.530 4.280 ;
        RECT 222.370 4.000 226.130 4.280 ;
        RECT 226.970 4.000 231.650 4.280 ;
        RECT 232.490 4.000 236.250 4.280 ;
        RECT 237.090 4.000 241.770 4.280 ;
        RECT 242.610 4.000 246.370 4.280 ;
        RECT 247.210 4.000 251.890 4.280 ;
        RECT 252.730 4.000 256.490 4.280 ;
        RECT 257.330 4.000 262.010 4.280 ;
        RECT 262.850 4.000 266.610 4.280 ;
        RECT 267.450 4.000 272.130 4.280 ;
        RECT 272.970 4.000 276.730 4.280 ;
        RECT 277.570 4.000 282.250 4.280 ;
        RECT 283.090 4.000 287.770 4.280 ;
        RECT 288.610 4.000 292.370 4.280 ;
        RECT 293.210 4.000 297.890 4.280 ;
        RECT 298.730 4.000 302.490 4.280 ;
        RECT 303.330 4.000 308.010 4.280 ;
        RECT 308.850 4.000 312.610 4.280 ;
        RECT 313.450 4.000 318.130 4.280 ;
        RECT 318.970 4.000 322.730 4.280 ;
        RECT 323.570 4.000 328.250 4.280 ;
        RECT 329.090 4.000 332.850 4.280 ;
        RECT 333.690 4.000 338.370 4.280 ;
        RECT 339.210 4.000 342.970 4.280 ;
        RECT 343.810 4.000 348.490 4.280 ;
        RECT 349.330 4.000 354.010 4.280 ;
        RECT 354.850 4.000 358.610 4.280 ;
        RECT 359.450 4.000 364.130 4.280 ;
        RECT 364.970 4.000 368.730 4.280 ;
        RECT 369.570 4.000 374.250 4.280 ;
        RECT 375.090 4.000 378.850 4.280 ;
        RECT 379.690 4.000 384.370 4.280 ;
        RECT 385.210 4.000 388.970 4.280 ;
        RECT 389.810 4.000 394.490 4.280 ;
        RECT 395.330 4.000 399.090 4.280 ;
        RECT 399.930 4.000 404.610 4.280 ;
        RECT 405.450 4.000 409.210 4.280 ;
        RECT 410.050 4.000 414.730 4.280 ;
        RECT 415.570 4.000 419.330 4.280 ;
        RECT 420.170 4.000 424.850 4.280 ;
        RECT 425.690 4.000 430.370 4.280 ;
        RECT 431.210 4.000 434.970 4.280 ;
        RECT 435.810 4.000 440.490 4.280 ;
        RECT 441.330 4.000 445.090 4.280 ;
        RECT 445.930 4.000 450.610 4.280 ;
        RECT 451.450 4.000 455.210 4.280 ;
        RECT 456.050 4.000 460.730 4.280 ;
        RECT 461.570 4.000 465.330 4.280 ;
        RECT 466.170 4.000 470.850 4.280 ;
        RECT 471.690 4.000 475.450 4.280 ;
        RECT 476.290 4.000 480.970 4.280 ;
        RECT 481.810 4.000 485.570 4.280 ;
        RECT 486.410 4.000 491.090 4.280 ;
        RECT 491.930 4.000 496.610 4.280 ;
      LAYER met3 ;
        RECT 3.990 505.560 495.550 506.425 ;
        RECT 3.990 501.520 495.950 505.560 ;
        RECT 4.400 500.160 495.950 501.520 ;
        RECT 4.400 500.120 495.550 500.160 ;
        RECT 3.990 498.760 495.550 500.120 ;
        RECT 3.990 493.360 495.950 498.760 ;
        RECT 4.400 492.000 495.950 493.360 ;
        RECT 4.400 491.960 495.550 492.000 ;
        RECT 3.990 490.600 495.550 491.960 ;
        RECT 3.990 486.560 495.950 490.600 ;
        RECT 4.400 485.200 495.950 486.560 ;
        RECT 4.400 485.160 495.550 485.200 ;
        RECT 3.990 483.800 495.550 485.160 ;
        RECT 3.990 478.400 495.950 483.800 ;
        RECT 4.400 477.040 495.950 478.400 ;
        RECT 4.400 477.000 495.550 477.040 ;
        RECT 3.990 475.640 495.550 477.000 ;
        RECT 3.990 471.600 495.950 475.640 ;
        RECT 4.400 470.240 495.950 471.600 ;
        RECT 4.400 470.200 495.550 470.240 ;
        RECT 3.990 468.840 495.550 470.200 ;
        RECT 3.990 463.440 495.950 468.840 ;
        RECT 4.400 462.080 495.950 463.440 ;
        RECT 4.400 462.040 495.550 462.080 ;
        RECT 3.990 460.680 495.550 462.040 ;
        RECT 3.990 456.640 495.950 460.680 ;
        RECT 4.400 455.280 495.950 456.640 ;
        RECT 4.400 455.240 495.550 455.280 ;
        RECT 3.990 453.880 495.550 455.240 ;
        RECT 3.990 448.480 495.950 453.880 ;
        RECT 4.400 447.120 495.950 448.480 ;
        RECT 4.400 447.080 495.550 447.120 ;
        RECT 3.990 445.720 495.550 447.080 ;
        RECT 3.990 441.680 495.950 445.720 ;
        RECT 4.400 440.320 495.950 441.680 ;
        RECT 4.400 440.280 495.550 440.320 ;
        RECT 3.990 438.920 495.550 440.280 ;
        RECT 3.990 433.520 495.950 438.920 ;
        RECT 4.400 432.160 495.950 433.520 ;
        RECT 4.400 432.120 495.550 432.160 ;
        RECT 3.990 430.760 495.550 432.120 ;
        RECT 3.990 426.720 495.950 430.760 ;
        RECT 4.400 425.360 495.950 426.720 ;
        RECT 4.400 425.320 495.550 425.360 ;
        RECT 3.990 423.960 495.550 425.320 ;
        RECT 3.990 418.560 495.950 423.960 ;
        RECT 4.400 417.200 495.950 418.560 ;
        RECT 4.400 417.160 495.550 417.200 ;
        RECT 3.990 415.800 495.550 417.160 ;
        RECT 3.990 410.400 495.950 415.800 ;
        RECT 4.400 409.000 495.550 410.400 ;
        RECT 3.990 403.600 495.950 409.000 ;
        RECT 4.400 402.240 495.950 403.600 ;
        RECT 4.400 402.200 495.550 402.240 ;
        RECT 3.990 400.840 495.550 402.200 ;
        RECT 3.990 395.440 495.950 400.840 ;
        RECT 4.400 394.080 495.950 395.440 ;
        RECT 4.400 394.040 495.550 394.080 ;
        RECT 3.990 392.680 495.550 394.040 ;
        RECT 3.990 388.640 495.950 392.680 ;
        RECT 4.400 387.280 495.950 388.640 ;
        RECT 4.400 387.240 495.550 387.280 ;
        RECT 3.990 385.880 495.550 387.240 ;
        RECT 3.990 380.480 495.950 385.880 ;
        RECT 4.400 379.120 495.950 380.480 ;
        RECT 4.400 379.080 495.550 379.120 ;
        RECT 3.990 377.720 495.550 379.080 ;
        RECT 3.990 373.680 495.950 377.720 ;
        RECT 4.400 372.320 495.950 373.680 ;
        RECT 4.400 372.280 495.550 372.320 ;
        RECT 3.990 370.920 495.550 372.280 ;
        RECT 3.990 365.520 495.950 370.920 ;
        RECT 4.400 364.160 495.950 365.520 ;
        RECT 4.400 364.120 495.550 364.160 ;
        RECT 3.990 362.760 495.550 364.120 ;
        RECT 3.990 358.720 495.950 362.760 ;
        RECT 4.400 357.360 495.950 358.720 ;
        RECT 4.400 357.320 495.550 357.360 ;
        RECT 3.990 355.960 495.550 357.320 ;
        RECT 3.990 350.560 495.950 355.960 ;
        RECT 4.400 349.200 495.950 350.560 ;
        RECT 4.400 349.160 495.550 349.200 ;
        RECT 3.990 347.800 495.550 349.160 ;
        RECT 3.990 343.760 495.950 347.800 ;
        RECT 4.400 342.400 495.950 343.760 ;
        RECT 4.400 342.360 495.550 342.400 ;
        RECT 3.990 341.000 495.550 342.360 ;
        RECT 3.990 335.600 495.950 341.000 ;
        RECT 4.400 334.240 495.950 335.600 ;
        RECT 4.400 334.200 495.550 334.240 ;
        RECT 3.990 332.840 495.550 334.200 ;
        RECT 3.990 328.800 495.950 332.840 ;
        RECT 4.400 327.440 495.950 328.800 ;
        RECT 4.400 327.400 495.550 327.440 ;
        RECT 3.990 326.040 495.550 327.400 ;
        RECT 3.990 320.640 495.950 326.040 ;
        RECT 4.400 319.280 495.950 320.640 ;
        RECT 4.400 319.240 495.550 319.280 ;
        RECT 3.990 317.880 495.550 319.240 ;
        RECT 3.990 313.840 495.950 317.880 ;
        RECT 4.400 312.480 495.950 313.840 ;
        RECT 4.400 312.440 495.550 312.480 ;
        RECT 3.990 311.080 495.550 312.440 ;
        RECT 3.990 305.680 495.950 311.080 ;
        RECT 4.400 304.320 495.950 305.680 ;
        RECT 4.400 304.280 495.550 304.320 ;
        RECT 3.990 302.920 495.550 304.280 ;
        RECT 3.990 297.520 495.950 302.920 ;
        RECT 4.400 296.160 495.950 297.520 ;
        RECT 4.400 296.120 495.550 296.160 ;
        RECT 3.990 294.760 495.550 296.120 ;
        RECT 3.990 290.720 495.950 294.760 ;
        RECT 4.400 289.360 495.950 290.720 ;
        RECT 4.400 289.320 495.550 289.360 ;
        RECT 3.990 287.960 495.550 289.320 ;
        RECT 3.990 282.560 495.950 287.960 ;
        RECT 4.400 281.200 495.950 282.560 ;
        RECT 4.400 281.160 495.550 281.200 ;
        RECT 3.990 279.800 495.550 281.160 ;
        RECT 3.990 275.760 495.950 279.800 ;
        RECT 4.400 274.400 495.950 275.760 ;
        RECT 4.400 274.360 495.550 274.400 ;
        RECT 3.990 273.000 495.550 274.360 ;
        RECT 3.990 267.600 495.950 273.000 ;
        RECT 4.400 266.240 495.950 267.600 ;
        RECT 4.400 266.200 495.550 266.240 ;
        RECT 3.990 264.840 495.550 266.200 ;
        RECT 3.990 260.800 495.950 264.840 ;
        RECT 4.400 259.440 495.950 260.800 ;
        RECT 4.400 259.400 495.550 259.440 ;
        RECT 3.990 258.040 495.550 259.400 ;
        RECT 3.990 252.640 495.950 258.040 ;
        RECT 4.400 251.280 495.950 252.640 ;
        RECT 4.400 251.240 495.550 251.280 ;
        RECT 3.990 249.880 495.550 251.240 ;
        RECT 3.990 245.840 495.950 249.880 ;
        RECT 4.400 244.480 495.950 245.840 ;
        RECT 4.400 244.440 495.550 244.480 ;
        RECT 3.990 243.080 495.550 244.440 ;
        RECT 3.990 237.680 495.950 243.080 ;
        RECT 4.400 236.320 495.950 237.680 ;
        RECT 4.400 236.280 495.550 236.320 ;
        RECT 3.990 234.920 495.550 236.280 ;
        RECT 3.990 230.880 495.950 234.920 ;
        RECT 4.400 229.520 495.950 230.880 ;
        RECT 4.400 229.480 495.550 229.520 ;
        RECT 3.990 228.120 495.550 229.480 ;
        RECT 3.990 222.720 495.950 228.120 ;
        RECT 4.400 221.360 495.950 222.720 ;
        RECT 4.400 221.320 495.550 221.360 ;
        RECT 3.990 219.960 495.550 221.320 ;
        RECT 3.990 215.920 495.950 219.960 ;
        RECT 4.400 214.560 495.950 215.920 ;
        RECT 4.400 214.520 495.550 214.560 ;
        RECT 3.990 213.160 495.550 214.520 ;
        RECT 3.990 207.760 495.950 213.160 ;
        RECT 4.400 206.400 495.950 207.760 ;
        RECT 4.400 206.360 495.550 206.400 ;
        RECT 3.990 205.000 495.550 206.360 ;
        RECT 3.990 199.600 495.950 205.000 ;
        RECT 4.400 198.200 495.550 199.600 ;
        RECT 3.990 192.800 495.950 198.200 ;
        RECT 4.400 191.440 495.950 192.800 ;
        RECT 4.400 191.400 495.550 191.440 ;
        RECT 3.990 190.040 495.550 191.400 ;
        RECT 3.990 184.640 495.950 190.040 ;
        RECT 4.400 183.280 495.950 184.640 ;
        RECT 4.400 183.240 495.550 183.280 ;
        RECT 3.990 181.880 495.550 183.240 ;
        RECT 3.990 177.840 495.950 181.880 ;
        RECT 4.400 176.480 495.950 177.840 ;
        RECT 4.400 176.440 495.550 176.480 ;
        RECT 3.990 175.080 495.550 176.440 ;
        RECT 3.990 169.680 495.950 175.080 ;
        RECT 4.400 168.320 495.950 169.680 ;
        RECT 4.400 168.280 495.550 168.320 ;
        RECT 3.990 166.920 495.550 168.280 ;
        RECT 3.990 162.880 495.950 166.920 ;
        RECT 4.400 161.520 495.950 162.880 ;
        RECT 4.400 161.480 495.550 161.520 ;
        RECT 3.990 160.120 495.550 161.480 ;
        RECT 3.990 154.720 495.950 160.120 ;
        RECT 4.400 153.360 495.950 154.720 ;
        RECT 4.400 153.320 495.550 153.360 ;
        RECT 3.990 151.960 495.550 153.320 ;
        RECT 3.990 147.920 495.950 151.960 ;
        RECT 4.400 146.560 495.950 147.920 ;
        RECT 4.400 146.520 495.550 146.560 ;
        RECT 3.990 145.160 495.550 146.520 ;
        RECT 3.990 139.760 495.950 145.160 ;
        RECT 4.400 138.400 495.950 139.760 ;
        RECT 4.400 138.360 495.550 138.400 ;
        RECT 3.990 137.000 495.550 138.360 ;
        RECT 3.990 132.960 495.950 137.000 ;
        RECT 4.400 131.600 495.950 132.960 ;
        RECT 4.400 131.560 495.550 131.600 ;
        RECT 3.990 130.200 495.550 131.560 ;
        RECT 3.990 124.800 495.950 130.200 ;
        RECT 4.400 123.440 495.950 124.800 ;
        RECT 4.400 123.400 495.550 123.440 ;
        RECT 3.990 122.040 495.550 123.400 ;
        RECT 3.990 118.000 495.950 122.040 ;
        RECT 4.400 116.640 495.950 118.000 ;
        RECT 4.400 116.600 495.550 116.640 ;
        RECT 3.990 115.240 495.550 116.600 ;
        RECT 3.990 109.840 495.950 115.240 ;
        RECT 4.400 108.480 495.950 109.840 ;
        RECT 4.400 108.440 495.550 108.480 ;
        RECT 3.990 107.080 495.550 108.440 ;
        RECT 3.990 101.680 495.950 107.080 ;
        RECT 4.400 100.280 495.550 101.680 ;
        RECT 3.990 94.880 495.950 100.280 ;
        RECT 4.400 93.520 495.950 94.880 ;
        RECT 4.400 93.480 495.550 93.520 ;
        RECT 3.990 92.120 495.550 93.480 ;
        RECT 3.990 86.720 495.950 92.120 ;
        RECT 4.400 85.360 495.950 86.720 ;
        RECT 4.400 85.320 495.550 85.360 ;
        RECT 3.990 83.960 495.550 85.320 ;
        RECT 3.990 79.920 495.950 83.960 ;
        RECT 4.400 78.560 495.950 79.920 ;
        RECT 4.400 78.520 495.550 78.560 ;
        RECT 3.990 77.160 495.550 78.520 ;
        RECT 3.990 71.760 495.950 77.160 ;
        RECT 4.400 70.400 495.950 71.760 ;
        RECT 4.400 70.360 495.550 70.400 ;
        RECT 3.990 69.000 495.550 70.360 ;
        RECT 3.990 64.960 495.950 69.000 ;
        RECT 4.400 63.600 495.950 64.960 ;
        RECT 4.400 63.560 495.550 63.600 ;
        RECT 3.990 62.200 495.550 63.560 ;
        RECT 3.990 56.800 495.950 62.200 ;
        RECT 4.400 55.440 495.950 56.800 ;
        RECT 4.400 55.400 495.550 55.440 ;
        RECT 3.990 54.040 495.550 55.400 ;
        RECT 3.990 50.000 495.950 54.040 ;
        RECT 4.400 48.640 495.950 50.000 ;
        RECT 4.400 48.600 495.550 48.640 ;
        RECT 3.990 47.240 495.550 48.600 ;
        RECT 3.990 41.840 495.950 47.240 ;
        RECT 4.400 40.480 495.950 41.840 ;
        RECT 4.400 40.440 495.550 40.480 ;
        RECT 3.990 39.080 495.550 40.440 ;
        RECT 3.990 35.040 495.950 39.080 ;
        RECT 4.400 33.680 495.950 35.040 ;
        RECT 4.400 33.640 495.550 33.680 ;
        RECT 3.990 32.280 495.550 33.640 ;
        RECT 3.990 26.880 495.950 32.280 ;
        RECT 4.400 25.520 495.950 26.880 ;
        RECT 4.400 25.480 495.550 25.520 ;
        RECT 3.990 24.120 495.550 25.480 ;
        RECT 3.990 20.080 495.950 24.120 ;
        RECT 4.400 18.720 495.950 20.080 ;
        RECT 4.400 18.680 495.550 18.720 ;
        RECT 3.990 17.320 495.550 18.680 ;
        RECT 3.990 11.920 495.950 17.320 ;
        RECT 4.400 10.560 495.950 11.920 ;
        RECT 4.400 10.520 495.550 10.560 ;
        RECT 3.990 9.160 495.550 10.520 ;
        RECT 3.990 4.255 495.950 9.160 ;
      LAYER met4 ;
        RECT 16.855 10.640 484.545 498.000 ;
      LAYER met5 ;
        RECT 5.520 106.280 494.040 487.630 ;
        RECT 5.520 29.690 494.040 101.480 ;
        RECT 5.520 17.900 494.040 24.890 ;
  END
END mac_cluster
END LIBRARY

