VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mac_cluster
  CLASS BLOCK ;
  FOREIGN mac_cluster ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.855 BY 511.575 ;
  PIN A0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.850 507.575 187.130 511.575 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 273.400 500.855 274.000 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 421.450 507.575 421.730 511.575 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.490 507.575 202.770 511.575 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END A0[7]
  PIN A1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.730 507.575 177.010 511.575 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 469.240 500.855 469.840 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.130 507.575 264.410 511.575 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.970 507.575 289.250 511.575 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 507.575 18.770 511.575 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.250 507.575 274.530 511.575 ;
    END
  END A1[7]
  PIN A2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 452.730 507.575 453.010 511.575 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END A2[6]
  PIN A2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 446.120 500.855 446.720 ;
    END
  END A2[7]
  PIN A3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 238.370 507.575 238.650 511.575 ;
    END
  END A3[0]
  PIN A3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END A3[1]
  PIN A3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 467.450 507.575 467.730 511.575 ;
    END
  END A3[2]
  PIN A3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.010 507.575 208.290 511.575 ;
    END
  END A3[3]
  PIN A3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END A3[4]
  PIN A3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END A3[5]
  PIN A3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END A3[6]
  PIN A3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.010 507.575 70.290 511.575 ;
    END
  END A3[7]
  PIN B0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END B0[0]
  PIN B0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END B0[1]
  PIN B0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END B0[2]
  PIN B0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END B0[3]
  PIN B0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 220.360 500.855 220.960 ;
    END
  END B0[4]
  PIN B0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.250 507.575 228.530 511.575 ;
    END
  END B0[5]
  PIN B0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 507.575 74.890 511.575 ;
    END
  END B0[6]
  PIN B0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END B0[7]
  PIN B1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 146.370 507.575 146.650 511.575 ;
    END
  END B1[0]
  PIN B1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 371.320 500.855 371.920 ;
    END
  END B1[1]
  PIN B1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 152.360 500.855 152.960 ;
    END
  END B1[2]
  PIN B1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END B1[3]
  PIN B1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 375.450 507.575 375.730 511.575 ;
    END
  END B1[4]
  PIN B1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END B1[5]
  PIN B1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.490 507.575 156.770 511.575 ;
    END
  END B1[6]
  PIN B1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 243.480 500.855 244.080 ;
    END
  END B1[7]
  PIN B2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END B2[0]
  PIN B2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END B2[1]
  PIN B2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END B2[2]
  PIN B2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 114.280 500.855 114.880 ;
    END
  END B2[3]
  PIN B2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 162.010 507.575 162.290 511.575 ;
    END
  END B2[4]
  PIN B2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 507.575 24.290 511.575 ;
    END
  END B2[5]
  PIN B2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END B2[6]
  PIN B2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 280.200 500.855 280.800 ;
    END
  END B2[7]
  PIN B3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 77.560 500.855 78.160 ;
    END
  END B3[0]
  PIN B3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END B3[1]
  PIN B3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END B3[2]
  PIN B3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 484.200 500.855 484.800 ;
    END
  END B3[3]
  PIN B3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 212.200 500.855 212.800 ;
    END
  END B3[4]
  PIN B3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 507.575 29.810 511.575 ;
    END
  END B3[5]
  PIN B3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END B3[6]
  PIN B3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 107.480 500.855 108.080 ;
    END
  END B3[7]
  PIN cfg[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.610 507.575 258.890 511.575 ;
    END
  END cfg[0]
  PIN cfg[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END cfg[100]
  PIN cfg[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END cfg[101]
  PIN cfg[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END cfg[102]
  PIN cfg[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 507.575 50.050 511.575 ;
    END
  END cfg[103]
  PIN cfg[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END cfg[104]
  PIN cfg[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END cfg[105]
  PIN cfg[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 431.160 500.855 431.760 ;
    END
  END cfg[106]
  PIN cfg[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END cfg[107]
  PIN cfg[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END cfg[108]
  PIN cfg[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 507.575 110.770 511.575 ;
    END
  END cfg[109]
  PIN cfg[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END cfg[10]
  PIN cfg[110]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END cfg[110]
  PIN cfg[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END cfg[111]
  PIN cfg[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END cfg[112]
  PIN cfg[113]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 205.400 500.855 206.000 ;
    END
  END cfg[113]
  PIN cfg[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 250.280 500.855 250.880 ;
    END
  END cfg[114]
  PIN cfg[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.250 507.575 90.530 511.575 ;
    END
  END cfg[115]
  PIN cfg[116]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END cfg[116]
  PIN cfg[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 431.570 507.575 431.850 511.575 ;
    END
  END cfg[117]
  PIN cfg[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END cfg[118]
  PIN cfg[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END cfg[119]
  PIN cfg[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END cfg[11]
  PIN cfg[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 120.610 507.575 120.890 511.575 ;
    END
  END cfg[120]
  PIN cfg[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 24.520 500.855 25.120 ;
    END
  END cfg[121]
  PIN cfg[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END cfg[122]
  PIN cfg[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END cfg[123]
  PIN cfg[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 363.160 500.855 363.760 ;
    END
  END cfg[124]
  PIN cfg[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 507.575 34.410 511.575 ;
    END
  END cfg[125]
  PIN cfg[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 258.440 500.855 259.040 ;
    END
  END cfg[126]
  PIN cfg[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END cfg[127]
  PIN cfg[128]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END cfg[128]
  PIN cfg[129]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END cfg[129]
  PIN cfg[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END cfg[12]
  PIN cfg[130]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END cfg[130]
  PIN cfg[131]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 350.610 507.575 350.890 511.575 ;
    END
  END cfg[131]
  PIN cfg[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 324.850 507.575 325.130 511.575 ;
    END
  END cfg[13]
  PIN cfg[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END cfg[14]
  PIN cfg[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END cfg[15]
  PIN cfg[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END cfg[16]
  PIN cfg[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 294.490 507.575 294.770 511.575 ;
    END
  END cfg[17]
  PIN cfg[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 356.360 500.855 356.960 ;
    END
  END cfg[18]
  PIN cfg[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END cfg[19]
  PIN cfg[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END cfg[1]
  PIN cfg[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 212.610 507.575 212.890 511.575 ;
    END
  END cfg[20]
  PIN cfg[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 92.520 500.855 93.120 ;
    END
  END cfg[21]
  PIN cfg[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 175.480 500.855 176.080 ;
    END
  END cfg[22]
  PIN cfg[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END cfg[23]
  PIN cfg[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 16.360 500.855 16.960 ;
    END
  END cfg[24]
  PIN cfg[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END cfg[25]
  PIN cfg[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END cfg[26]
  PIN cfg[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 340.490 507.575 340.770 511.575 ;
    END
  END cfg[27]
  PIN cfg[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 437.090 507.575 437.370 511.575 ;
    END
  END cfg[28]
  PIN cfg[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END cfg[29]
  PIN cfg[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END cfg[2]
  PIN cfg[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END cfg[30]
  PIN cfg[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 318.280 500.855 318.880 ;
    END
  END cfg[31]
  PIN cfg[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.970 507.575 473.250 511.575 ;
    END
  END cfg[32]
  PIN cfg[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 253.090 507.575 253.370 511.575 ;
    END
  END cfg[33]
  PIN cfg[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END cfg[34]
  PIN cfg[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END cfg[35]
  PIN cfg[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END cfg[36]
  PIN cfg[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END cfg[37]
  PIN cfg[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 54.440 500.855 55.040 ;
    END
  END cfg[38]
  PIN cfg[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 386.280 500.855 386.880 ;
    END
  END cfg[39]
  PIN cfg[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 461.080 500.855 461.680 ;
    END
  END cfg[3]
  PIN cfg[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END cfg[40]
  PIN cfg[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 507.575 85.930 511.575 ;
    END
  END cfg[41]
  PIN cfg[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END cfg[42]
  PIN cfg[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END cfg[43]
  PIN cfg[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 129.240 500.855 129.840 ;
    END
  END cfg[44]
  PIN cfg[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END cfg[45]
  PIN cfg[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 408.040 500.855 408.640 ;
    END
  END cfg[46]
  PIN cfg[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.210 507.575 401.490 511.575 ;
    END
  END cfg[47]
  PIN cfg[48]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END cfg[48]
  PIN cfg[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 507.575 80.410 511.575 ;
    END
  END cfg[49]
  PIN cfg[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.130 507.575 172.410 511.575 ;
    END
  END cfg[4]
  PIN cfg[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END cfg[50]
  PIN cfg[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.850 507.575 463.130 511.575 ;
    END
  END cfg[51]
  PIN cfg[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END cfg[52]
  PIN cfg[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END cfg[53]
  PIN cfg[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END cfg[54]
  PIN cfg[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END cfg[55]
  PIN cfg[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END cfg[56]
  PIN cfg[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END cfg[57]
  PIN cfg[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.490 507.575 386.770 511.575 ;
    END
  END cfg[58]
  PIN cfg[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END cfg[59]
  PIN cfg[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 391.090 507.575 391.370 511.575 ;
    END
  END cfg[5]
  PIN cfg[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 491.000 500.855 491.600 ;
    END
  END cfg[60]
  PIN cfg[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 295.160 500.855 295.760 ;
    END
  END cfg[61]
  PIN cfg[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.090 507.575 299.370 511.575 ;
    END
  END cfg[62]
  PIN cfg[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 144.200 500.855 144.800 ;
    END
  END cfg[63]
  PIN cfg[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END cfg[64]
  PIN cfg[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END cfg[65]
  PIN cfg[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 507.575 106.170 511.575 ;
    END
  END cfg[66]
  PIN cfg[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 507.575 4.050 511.575 ;
    END
  END cfg[67]
  PIN cfg[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END cfg[68]
  PIN cfg[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END cfg[69]
  PIN cfg[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 304.610 507.575 304.890 511.575 ;
    END
  END cfg[6]
  PIN cfg[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END cfg[70]
  PIN cfg[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 160.520 500.855 161.120 ;
    END
  END cfg[71]
  PIN cfg[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END cfg[72]
  PIN cfg[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END cfg[73]
  PIN cfg[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.610 507.575 166.890 511.575 ;
    END
  END cfg[74]
  PIN cfg[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END cfg[75]
  PIN cfg[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END cfg[76]
  PIN cfg[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END cfg[77]
  PIN cfg[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 31.320 500.855 31.920 ;
    END
  END cfg[78]
  PIN cfg[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 406.730 507.575 407.010 511.575 ;
    END
  END cfg[79]
  PIN cfg[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END cfg[7]
  PIN cfg[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END cfg[80]
  PIN cfg[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END cfg[81]
  PIN cfg[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END cfg[82]
  PIN cfg[83]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END cfg[83]
  PIN cfg[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 497.810 507.575 498.090 511.575 ;
    END
  END cfg[84]
  PIN cfg[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 360.730 507.575 361.010 511.575 ;
    END
  END cfg[85]
  PIN cfg[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 320.250 507.575 320.530 511.575 ;
    END
  END cfg[86]
  PIN cfg[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 197.240 500.855 197.840 ;
    END
  END cfg[87]
  PIN cfg[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.970 507.575 335.250 511.575 ;
    END
  END cfg[88]
  PIN cfg[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END cfg[89]
  PIN cfg[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 333.240 500.855 333.840 ;
    END
  END cfg[8]
  PIN cfg[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END cfg[90]
  PIN cfg[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END cfg[91]
  PIN cfg[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END cfg[92]
  PIN cfg[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END cfg[93]
  PIN cfg[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END cfg[94]
  PIN cfg[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.010 507.575 116.290 511.575 ;
    END
  END cfg[95]
  PIN cfg[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 99.320 500.855 99.920 ;
    END
  END cfg[96]
  PIN cfg[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END cfg[97]
  PIN cfg[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END cfg[98]
  PIN cfg[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END cfg[99]
  PIN cfg[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 416.200 500.855 416.800 ;
    END
  END cfg[9]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.570 507.575 477.850 511.575 ;
    END
  END clk
  PIN cset
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 496.855 227.160 500.855 227.760 ;
    END
  END cset
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 278.850 507.575 279.130 511.575 ;
    END
  END en
  PIN out0[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END out0[0]
  PIN out0[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 416.850 507.575 417.130 511.575 ;
    END
  END out0[10]
  PIN out0[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 265.240 500.855 265.840 ;
    END
  END out0[11]
  PIN out0[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 424.360 500.855 424.960 ;
    END
  END out0[12]
  PIN out0[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 303.320 500.855 303.920 ;
    END
  END out0[13]
  PIN out0[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 122.440 500.855 123.040 ;
    END
  END out0[14]
  PIN out0[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 182.250 507.575 182.530 511.575 ;
    END
  END out0[15]
  PIN out0[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 141.770 507.575 142.050 511.575 ;
    END
  END out0[16]
  PIN out0[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.130 507.575 126.410 511.575 ;
    END
  END out0[17]
  PIN out0[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END out0[18]
  PIN out0[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 415.010 0.000 415.290 4.000 ;
    END
  END out0[19]
  PIN out0[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 341.400 500.855 342.000 ;
    END
  END out0[1]
  PIN out0[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END out0[20]
  PIN out0[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END out0[21]
  PIN out0[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END out0[22]
  PIN out0[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END out0[23]
  PIN out0[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.730 507.575 223.010 511.575 ;
    END
  END out0[24]
  PIN out0[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 380.970 507.575 381.250 511.575 ;
    END
  END out0[25]
  PIN out0[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 401.240 500.855 401.840 ;
    END
  END out0[26]
  PIN out0[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 454.280 500.855 454.880 ;
    END
  END out0[27]
  PIN out0[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.370 507.575 54.650 511.575 ;
    END
  END out0[28]
  PIN out0[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 325.080 500.855 325.680 ;
    END
  END out0[29]
  PIN out0[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 457.330 507.575 457.610 511.575 ;
    END
  END out0[2]
  PIN out0[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END out0[30]
  PIN out0[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END out0[31]
  PIN out0[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END out0[3]
  PIN out0[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 39.480 500.855 40.080 ;
    END
  END out0[4]
  PIN out0[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 378.120 500.855 378.720 ;
    END
  END out0[5]
  PIN out0[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 345.090 507.575 345.370 511.575 ;
    END
  END out0[6]
  PIN out0[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 310.120 500.855 310.720 ;
    END
  END out0[7]
  PIN out0[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END out0[8]
  PIN out0[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 487.690 507.575 487.970 511.575 ;
    END
  END out0[9]
  PIN out1[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 330.370 507.575 330.650 511.575 ;
    END
  END out1[0]
  PIN out1[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 348.200 500.855 348.800 ;
    END
  END out1[10]
  PIN out1[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 439.320 500.855 439.920 ;
    END
  END out1[11]
  PIN out1[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END out1[12]
  PIN out1[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END out1[13]
  PIN out1[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.250 507.575 44.530 511.575 ;
    END
  END out1[14]
  PIN out1[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 309.210 507.575 309.490 511.575 ;
    END
  END out1[15]
  PIN out1[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END out1[16]
  PIN out1[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 190.440 500.855 191.040 ;
    END
  END out1[17]
  PIN out1[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.650 507.575 39.930 511.575 ;
    END
  END out1[18]
  PIN out1[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END out1[19]
  PIN out1[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END out1[1]
  PIN out1[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 476.040 500.855 476.640 ;
    END
  END out1[20]
  PIN out1[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 426.970 507.575 427.250 511.575 ;
    END
  END out1[21]
  PIN out1[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END out1[22]
  PIN out1[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END out1[23]
  PIN out1[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 507.575 131.010 511.575 ;
    END
  END out1[24]
  PIN out1[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END out1[25]
  PIN out1[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END out1[26]
  PIN out1[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 483.090 507.575 483.370 511.575 ;
    END
  END out1[27]
  PIN out1[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 167.320 500.855 167.920 ;
    END
  END out1[28]
  PIN out1[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END out1[29]
  PIN out1[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END out1[2]
  PIN out1[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END out1[30]
  PIN out1[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 507.575 14.170 511.575 ;
    END
  END out1[31]
  PIN out1[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 69.400 500.855 70.000 ;
    END
  END out1[3]
  PIN out1[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END out1[4]
  PIN out1[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END out1[5]
  PIN out1[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END out1[6]
  PIN out1[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 182.280 500.855 182.880 ;
    END
  END out1[7]
  PIN out1[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 218.130 507.575 218.410 511.575 ;
    END
  END out1[8]
  PIN out1[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.250 507.575 136.530 511.575 ;
    END
  END out1[9]
  PIN out2[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END out2[0]
  PIN out2[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END out2[10]
  PIN out2[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 507.575 100.650 511.575 ;
    END
  END out2[11]
  PIN out2[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 137.400 500.855 138.000 ;
    END
  END out2[12]
  PIN out2[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END out2[13]
  PIN out2[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END out2[14]
  PIN out2[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 248.490 507.575 248.770 511.575 ;
    END
  END out2[15]
  PIN out2[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 314.730 507.575 315.010 511.575 ;
    END
  END out2[16]
  PIN out2[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END out2[17]
  PIN out2[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 393.080 500.855 393.680 ;
    END
  END out2[18]
  PIN out2[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END out2[19]
  PIN out2[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END out2[1]
  PIN out2[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 151.890 507.575 152.170 511.575 ;
    END
  END out2[20]
  PIN out2[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END out2[21]
  PIN out2[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 499.160 500.855 499.760 ;
    END
  END out2[22]
  PIN out2[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END out2[23]
  PIN out2[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 235.320 500.855 235.920 ;
    END
  END out2[24]
  PIN out2[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END out2[25]
  PIN out2[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 46.280 500.855 46.880 ;
    END
  END out2[26]
  PIN out2[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END out2[27]
  PIN out2[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 447.210 507.575 447.490 511.575 ;
    END
  END out2[28]
  PIN out2[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END out2[29]
  PIN out2[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 242.970 507.575 243.250 511.575 ;
    END
  END out2[2]
  PIN out2[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END out2[30]
  PIN out2[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END out2[31]
  PIN out2[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.490 507.575 64.770 511.575 ;
    END
  END out2[3]
  PIN out2[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 396.610 507.575 396.890 511.575 ;
    END
  END out2[4]
  PIN out2[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 192.370 507.575 192.650 511.575 ;
    END
  END out2[5]
  PIN out2[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END out2[6]
  PIN out2[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.970 507.575 197.250 511.575 ;
    END
  END out2[7]
  PIN out2[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END out2[8]
  PIN out2[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 61.240 500.855 61.840 ;
    END
  END out2[9]
  PIN out3[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END out3[0]
  PIN out3[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 442.610 507.575 442.890 511.575 ;
    END
  END out3[10]
  PIN out3[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 284.370 507.575 284.650 511.575 ;
    END
  END out3[11]
  PIN out3[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 355.210 507.575 355.490 511.575 ;
    END
  END out3[12]
  PIN out3[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END out3[13]
  PIN out3[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END out3[14]
  PIN out3[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 288.360 500.855 288.960 ;
    END
  END out3[15]
  PIN out3[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END out3[16]
  PIN out3[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END out3[17]
  PIN out3[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 365.330 507.575 365.610 511.575 ;
    END
  END out3[18]
  PIN out3[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 507.575 96.050 511.575 ;
    END
  END out3[19]
  PIN out3[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 507.575 60.170 511.575 ;
    END
  END out3[1]
  PIN out3[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END out3[20]
  PIN out3[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END out3[21]
  PIN out3[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END out3[22]
  PIN out3[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 268.730 507.575 269.010 511.575 ;
    END
  END out3[23]
  PIN out3[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END out3[24]
  PIN out3[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 84.360 500.855 84.960 ;
    END
  END out3[25]
  PIN out3[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END out3[26]
  PIN out3[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 507.575 8.650 511.575 ;
    END
  END out3[27]
  PIN out3[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 370.850 507.575 371.130 511.575 ;
    END
  END out3[28]
  PIN out3[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 411.330 507.575 411.610 511.575 ;
    END
  END out3[29]
  PIN out3[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END out3[2]
  PIN out3[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END out3[30]
  PIN out3[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END out3[31]
  PIN out3[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END out3[3]
  PIN out3[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END out3[4]
  PIN out3[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 232.850 507.575 233.130 511.575 ;
    END
  END out3[5]
  PIN out3[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END out3[6]
  PIN out3[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 496.855 9.560 500.855 10.160 ;
    END
  END out3[7]
  PIN out3[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END out3[8]
  PIN out3[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 493.210 507.575 493.490 511.575 ;
    END
  END out3[9]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END rst
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 494.960 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 494.960 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.960 500.565 ;
      LAYER met1 ;
        RECT 0.530 6.160 498.110 507.240 ;
      LAYER met2 ;
        RECT 0.160 507.295 3.490 507.575 ;
        RECT 4.330 507.295 8.090 507.575 ;
        RECT 8.930 507.295 13.610 507.575 ;
        RECT 14.450 507.295 18.210 507.575 ;
        RECT 19.050 507.295 23.730 507.575 ;
        RECT 24.570 507.295 29.250 507.575 ;
        RECT 30.090 507.295 33.850 507.575 ;
        RECT 34.690 507.295 39.370 507.575 ;
        RECT 40.210 507.295 43.970 507.575 ;
        RECT 44.810 507.295 49.490 507.575 ;
        RECT 50.330 507.295 54.090 507.575 ;
        RECT 54.930 507.295 59.610 507.575 ;
        RECT 60.450 507.295 64.210 507.575 ;
        RECT 65.050 507.295 69.730 507.575 ;
        RECT 70.570 507.295 74.330 507.575 ;
        RECT 75.170 507.295 79.850 507.575 ;
        RECT 80.690 507.295 85.370 507.575 ;
        RECT 86.210 507.295 89.970 507.575 ;
        RECT 90.810 507.295 95.490 507.575 ;
        RECT 96.330 507.295 100.090 507.575 ;
        RECT 100.930 507.295 105.610 507.575 ;
        RECT 106.450 507.295 110.210 507.575 ;
        RECT 111.050 507.295 115.730 507.575 ;
        RECT 116.570 507.295 120.330 507.575 ;
        RECT 121.170 507.295 125.850 507.575 ;
        RECT 126.690 507.295 130.450 507.575 ;
        RECT 131.290 507.295 135.970 507.575 ;
        RECT 136.810 507.295 141.490 507.575 ;
        RECT 142.330 507.295 146.090 507.575 ;
        RECT 146.930 507.295 151.610 507.575 ;
        RECT 152.450 507.295 156.210 507.575 ;
        RECT 157.050 507.295 161.730 507.575 ;
        RECT 162.570 507.295 166.330 507.575 ;
        RECT 167.170 507.295 171.850 507.575 ;
        RECT 172.690 507.295 176.450 507.575 ;
        RECT 177.290 507.295 181.970 507.575 ;
        RECT 182.810 507.295 186.570 507.575 ;
        RECT 187.410 507.295 192.090 507.575 ;
        RECT 192.930 507.295 196.690 507.575 ;
        RECT 197.530 507.295 202.210 507.575 ;
        RECT 203.050 507.295 207.730 507.575 ;
        RECT 208.570 507.295 212.330 507.575 ;
        RECT 213.170 507.295 217.850 507.575 ;
        RECT 218.690 507.295 222.450 507.575 ;
        RECT 223.290 507.295 227.970 507.575 ;
        RECT 228.810 507.295 232.570 507.575 ;
        RECT 233.410 507.295 238.090 507.575 ;
        RECT 238.930 507.295 242.690 507.575 ;
        RECT 243.530 507.295 248.210 507.575 ;
        RECT 249.050 507.295 252.810 507.575 ;
        RECT 253.650 507.295 258.330 507.575 ;
        RECT 259.170 507.295 263.850 507.575 ;
        RECT 264.690 507.295 268.450 507.575 ;
        RECT 269.290 507.295 273.970 507.575 ;
        RECT 274.810 507.295 278.570 507.575 ;
        RECT 279.410 507.295 284.090 507.575 ;
        RECT 284.930 507.295 288.690 507.575 ;
        RECT 289.530 507.295 294.210 507.575 ;
        RECT 295.050 507.295 298.810 507.575 ;
        RECT 299.650 507.295 304.330 507.575 ;
        RECT 305.170 507.295 308.930 507.575 ;
        RECT 309.770 507.295 314.450 507.575 ;
        RECT 315.290 507.295 319.970 507.575 ;
        RECT 320.810 507.295 324.570 507.575 ;
        RECT 325.410 507.295 330.090 507.575 ;
        RECT 330.930 507.295 334.690 507.575 ;
        RECT 335.530 507.295 340.210 507.575 ;
        RECT 341.050 507.295 344.810 507.575 ;
        RECT 345.650 507.295 350.330 507.575 ;
        RECT 351.170 507.295 354.930 507.575 ;
        RECT 355.770 507.295 360.450 507.575 ;
        RECT 361.290 507.295 365.050 507.575 ;
        RECT 365.890 507.295 370.570 507.575 ;
        RECT 371.410 507.295 375.170 507.575 ;
        RECT 376.010 507.295 380.690 507.575 ;
        RECT 381.530 507.295 386.210 507.575 ;
        RECT 387.050 507.295 390.810 507.575 ;
        RECT 391.650 507.295 396.330 507.575 ;
        RECT 397.170 507.295 400.930 507.575 ;
        RECT 401.770 507.295 406.450 507.575 ;
        RECT 407.290 507.295 411.050 507.575 ;
        RECT 411.890 507.295 416.570 507.575 ;
        RECT 417.410 507.295 421.170 507.575 ;
        RECT 422.010 507.295 426.690 507.575 ;
        RECT 427.530 507.295 431.290 507.575 ;
        RECT 432.130 507.295 436.810 507.575 ;
        RECT 437.650 507.295 442.330 507.575 ;
        RECT 443.170 507.295 446.930 507.575 ;
        RECT 447.770 507.295 452.450 507.575 ;
        RECT 453.290 507.295 457.050 507.575 ;
        RECT 457.890 507.295 462.570 507.575 ;
        RECT 463.410 507.295 467.170 507.575 ;
        RECT 468.010 507.295 472.690 507.575 ;
        RECT 473.530 507.295 477.290 507.575 ;
        RECT 478.130 507.295 482.810 507.575 ;
        RECT 483.650 507.295 487.410 507.575 ;
        RECT 488.250 507.295 492.930 507.575 ;
        RECT 493.770 507.295 497.530 507.575 ;
        RECT 0.160 4.280 498.080 507.295 ;
        RECT 0.160 4.000 2.570 4.280 ;
        RECT 3.410 4.000 7.170 4.280 ;
        RECT 8.010 4.000 12.690 4.280 ;
        RECT 13.530 4.000 17.290 4.280 ;
        RECT 18.130 4.000 22.810 4.280 ;
        RECT 23.650 4.000 27.410 4.280 ;
        RECT 28.250 4.000 32.930 4.280 ;
        RECT 33.770 4.000 37.530 4.280 ;
        RECT 38.370 4.000 43.050 4.280 ;
        RECT 43.890 4.000 47.650 4.280 ;
        RECT 48.490 4.000 53.170 4.280 ;
        RECT 54.010 4.000 57.770 4.280 ;
        RECT 58.610 4.000 63.290 4.280 ;
        RECT 64.130 4.000 68.810 4.280 ;
        RECT 69.650 4.000 73.410 4.280 ;
        RECT 74.250 4.000 78.930 4.280 ;
        RECT 79.770 4.000 83.530 4.280 ;
        RECT 84.370 4.000 89.050 4.280 ;
        RECT 89.890 4.000 93.650 4.280 ;
        RECT 94.490 4.000 99.170 4.280 ;
        RECT 100.010 4.000 103.770 4.280 ;
        RECT 104.610 4.000 109.290 4.280 ;
        RECT 110.130 4.000 113.890 4.280 ;
        RECT 114.730 4.000 119.410 4.280 ;
        RECT 120.250 4.000 124.930 4.280 ;
        RECT 125.770 4.000 129.530 4.280 ;
        RECT 130.370 4.000 135.050 4.280 ;
        RECT 135.890 4.000 139.650 4.280 ;
        RECT 140.490 4.000 145.170 4.280 ;
        RECT 146.010 4.000 149.770 4.280 ;
        RECT 150.610 4.000 155.290 4.280 ;
        RECT 156.130 4.000 159.890 4.280 ;
        RECT 160.730 4.000 165.410 4.280 ;
        RECT 166.250 4.000 170.010 4.280 ;
        RECT 170.850 4.000 175.530 4.280 ;
        RECT 176.370 4.000 180.130 4.280 ;
        RECT 180.970 4.000 185.650 4.280 ;
        RECT 186.490 4.000 191.170 4.280 ;
        RECT 192.010 4.000 195.770 4.280 ;
        RECT 196.610 4.000 201.290 4.280 ;
        RECT 202.130 4.000 205.890 4.280 ;
        RECT 206.730 4.000 211.410 4.280 ;
        RECT 212.250 4.000 216.010 4.280 ;
        RECT 216.850 4.000 221.530 4.280 ;
        RECT 222.370 4.000 226.130 4.280 ;
        RECT 226.970 4.000 231.650 4.280 ;
        RECT 232.490 4.000 236.250 4.280 ;
        RECT 237.090 4.000 241.770 4.280 ;
        RECT 242.610 4.000 247.290 4.280 ;
        RECT 248.130 4.000 251.890 4.280 ;
        RECT 252.730 4.000 257.410 4.280 ;
        RECT 258.250 4.000 262.010 4.280 ;
        RECT 262.850 4.000 267.530 4.280 ;
        RECT 268.370 4.000 272.130 4.280 ;
        RECT 272.970 4.000 277.650 4.280 ;
        RECT 278.490 4.000 282.250 4.280 ;
        RECT 283.090 4.000 287.770 4.280 ;
        RECT 288.610 4.000 292.370 4.280 ;
        RECT 293.210 4.000 297.890 4.280 ;
        RECT 298.730 4.000 303.410 4.280 ;
        RECT 304.250 4.000 308.010 4.280 ;
        RECT 308.850 4.000 313.530 4.280 ;
        RECT 314.370 4.000 318.130 4.280 ;
        RECT 318.970 4.000 323.650 4.280 ;
        RECT 324.490 4.000 328.250 4.280 ;
        RECT 329.090 4.000 333.770 4.280 ;
        RECT 334.610 4.000 338.370 4.280 ;
        RECT 339.210 4.000 343.890 4.280 ;
        RECT 344.730 4.000 348.490 4.280 ;
        RECT 349.330 4.000 354.010 4.280 ;
        RECT 354.850 4.000 358.610 4.280 ;
        RECT 359.450 4.000 364.130 4.280 ;
        RECT 364.970 4.000 369.650 4.280 ;
        RECT 370.490 4.000 374.250 4.280 ;
        RECT 375.090 4.000 379.770 4.280 ;
        RECT 380.610 4.000 384.370 4.280 ;
        RECT 385.210 4.000 389.890 4.280 ;
        RECT 390.730 4.000 394.490 4.280 ;
        RECT 395.330 4.000 400.010 4.280 ;
        RECT 400.850 4.000 404.610 4.280 ;
        RECT 405.450 4.000 410.130 4.280 ;
        RECT 410.970 4.000 414.730 4.280 ;
        RECT 415.570 4.000 420.250 4.280 ;
        RECT 421.090 4.000 425.770 4.280 ;
        RECT 426.610 4.000 430.370 4.280 ;
        RECT 431.210 4.000 435.890 4.280 ;
        RECT 436.730 4.000 440.490 4.280 ;
        RECT 441.330 4.000 446.010 4.280 ;
        RECT 446.850 4.000 450.610 4.280 ;
        RECT 451.450 4.000 456.130 4.280 ;
        RECT 456.970 4.000 460.730 4.280 ;
        RECT 461.570 4.000 466.250 4.280 ;
        RECT 467.090 4.000 470.850 4.280 ;
        RECT 471.690 4.000 476.370 4.280 ;
        RECT 477.210 4.000 481.890 4.280 ;
        RECT 482.730 4.000 486.490 4.280 ;
        RECT 487.330 4.000 492.010 4.280 ;
        RECT 492.850 4.000 496.610 4.280 ;
        RECT 497.450 4.000 498.080 4.280 ;
      LAYER met3 ;
        RECT 4.400 500.160 496.855 500.985 ;
        RECT 4.400 500.120 496.455 500.160 ;
        RECT 0.310 498.760 496.455 500.120 ;
        RECT 0.310 494.720 496.855 498.760 ;
        RECT 4.400 493.320 496.855 494.720 ;
        RECT 0.310 492.000 496.855 493.320 ;
        RECT 0.310 490.600 496.455 492.000 ;
        RECT 0.310 486.560 496.855 490.600 ;
        RECT 4.400 485.200 496.855 486.560 ;
        RECT 4.400 485.160 496.455 485.200 ;
        RECT 0.310 483.800 496.455 485.160 ;
        RECT 0.310 479.760 496.855 483.800 ;
        RECT 4.400 478.360 496.855 479.760 ;
        RECT 0.310 477.040 496.855 478.360 ;
        RECT 0.310 475.640 496.455 477.040 ;
        RECT 0.310 471.600 496.855 475.640 ;
        RECT 4.400 470.240 496.855 471.600 ;
        RECT 4.400 470.200 496.455 470.240 ;
        RECT 0.310 468.840 496.455 470.200 ;
        RECT 0.310 464.800 496.855 468.840 ;
        RECT 4.400 463.400 496.855 464.800 ;
        RECT 0.310 462.080 496.855 463.400 ;
        RECT 0.310 460.680 496.455 462.080 ;
        RECT 0.310 456.640 496.855 460.680 ;
        RECT 4.400 455.280 496.855 456.640 ;
        RECT 4.400 455.240 496.455 455.280 ;
        RECT 0.310 453.880 496.455 455.240 ;
        RECT 0.310 449.840 496.855 453.880 ;
        RECT 4.400 448.440 496.855 449.840 ;
        RECT 0.310 447.120 496.855 448.440 ;
        RECT 0.310 445.720 496.455 447.120 ;
        RECT 0.310 441.680 496.855 445.720 ;
        RECT 4.400 440.320 496.855 441.680 ;
        RECT 4.400 440.280 496.455 440.320 ;
        RECT 0.310 438.920 496.455 440.280 ;
        RECT 0.310 433.520 496.855 438.920 ;
        RECT 4.400 432.160 496.855 433.520 ;
        RECT 4.400 432.120 496.455 432.160 ;
        RECT 0.310 430.760 496.455 432.120 ;
        RECT 0.310 426.720 496.855 430.760 ;
        RECT 4.400 425.360 496.855 426.720 ;
        RECT 4.400 425.320 496.455 425.360 ;
        RECT 0.310 423.960 496.455 425.320 ;
        RECT 0.310 418.560 496.855 423.960 ;
        RECT 4.400 417.200 496.855 418.560 ;
        RECT 4.400 417.160 496.455 417.200 ;
        RECT 0.310 415.800 496.455 417.160 ;
        RECT 0.310 411.760 496.855 415.800 ;
        RECT 4.400 410.360 496.855 411.760 ;
        RECT 0.310 409.040 496.855 410.360 ;
        RECT 0.310 407.640 496.455 409.040 ;
        RECT 0.310 403.600 496.855 407.640 ;
        RECT 4.400 402.240 496.855 403.600 ;
        RECT 4.400 402.200 496.455 402.240 ;
        RECT 0.310 400.840 496.455 402.200 ;
        RECT 0.310 396.800 496.855 400.840 ;
        RECT 4.400 395.400 496.855 396.800 ;
        RECT 0.310 394.080 496.855 395.400 ;
        RECT 0.310 392.680 496.455 394.080 ;
        RECT 0.310 388.640 496.855 392.680 ;
        RECT 4.400 387.280 496.855 388.640 ;
        RECT 4.400 387.240 496.455 387.280 ;
        RECT 0.310 385.880 496.455 387.240 ;
        RECT 0.310 381.840 496.855 385.880 ;
        RECT 4.400 380.440 496.855 381.840 ;
        RECT 0.310 379.120 496.855 380.440 ;
        RECT 0.310 377.720 496.455 379.120 ;
        RECT 0.310 373.680 496.855 377.720 ;
        RECT 4.400 372.320 496.855 373.680 ;
        RECT 4.400 372.280 496.455 372.320 ;
        RECT 0.310 370.920 496.455 372.280 ;
        RECT 0.310 366.880 496.855 370.920 ;
        RECT 4.400 365.480 496.855 366.880 ;
        RECT 0.310 364.160 496.855 365.480 ;
        RECT 0.310 362.760 496.455 364.160 ;
        RECT 0.310 358.720 496.855 362.760 ;
        RECT 4.400 357.360 496.855 358.720 ;
        RECT 4.400 357.320 496.455 357.360 ;
        RECT 0.310 355.960 496.455 357.320 ;
        RECT 0.310 350.560 496.855 355.960 ;
        RECT 4.400 349.200 496.855 350.560 ;
        RECT 4.400 349.160 496.455 349.200 ;
        RECT 0.310 347.800 496.455 349.160 ;
        RECT 0.310 343.760 496.855 347.800 ;
        RECT 4.400 342.400 496.855 343.760 ;
        RECT 4.400 342.360 496.455 342.400 ;
        RECT 0.310 341.000 496.455 342.360 ;
        RECT 0.310 335.600 496.855 341.000 ;
        RECT 4.400 334.240 496.855 335.600 ;
        RECT 4.400 334.200 496.455 334.240 ;
        RECT 0.310 332.840 496.455 334.200 ;
        RECT 0.310 328.800 496.855 332.840 ;
        RECT 4.400 327.400 496.855 328.800 ;
        RECT 0.310 326.080 496.855 327.400 ;
        RECT 0.310 324.680 496.455 326.080 ;
        RECT 0.310 320.640 496.855 324.680 ;
        RECT 4.400 319.280 496.855 320.640 ;
        RECT 4.400 319.240 496.455 319.280 ;
        RECT 0.310 317.880 496.455 319.240 ;
        RECT 0.310 313.840 496.855 317.880 ;
        RECT 4.400 312.440 496.855 313.840 ;
        RECT 0.310 311.120 496.855 312.440 ;
        RECT 0.310 309.720 496.455 311.120 ;
        RECT 0.310 305.680 496.855 309.720 ;
        RECT 4.400 304.320 496.855 305.680 ;
        RECT 4.400 304.280 496.455 304.320 ;
        RECT 0.310 302.920 496.455 304.280 ;
        RECT 0.310 298.880 496.855 302.920 ;
        RECT 4.400 297.480 496.855 298.880 ;
        RECT 0.310 296.160 496.855 297.480 ;
        RECT 0.310 294.760 496.455 296.160 ;
        RECT 0.310 290.720 496.855 294.760 ;
        RECT 4.400 289.360 496.855 290.720 ;
        RECT 4.400 289.320 496.455 289.360 ;
        RECT 0.310 287.960 496.455 289.320 ;
        RECT 0.310 283.920 496.855 287.960 ;
        RECT 4.400 282.520 496.855 283.920 ;
        RECT 0.310 281.200 496.855 282.520 ;
        RECT 0.310 279.800 496.455 281.200 ;
        RECT 0.310 275.760 496.855 279.800 ;
        RECT 4.400 274.400 496.855 275.760 ;
        RECT 4.400 274.360 496.455 274.400 ;
        RECT 0.310 273.000 496.455 274.360 ;
        RECT 0.310 267.600 496.855 273.000 ;
        RECT 4.400 266.240 496.855 267.600 ;
        RECT 4.400 266.200 496.455 266.240 ;
        RECT 0.310 264.840 496.455 266.200 ;
        RECT 0.310 260.800 496.855 264.840 ;
        RECT 4.400 259.440 496.855 260.800 ;
        RECT 4.400 259.400 496.455 259.440 ;
        RECT 0.310 258.040 496.455 259.400 ;
        RECT 0.310 252.640 496.855 258.040 ;
        RECT 4.400 251.280 496.855 252.640 ;
        RECT 4.400 251.240 496.455 251.280 ;
        RECT 0.310 249.880 496.455 251.240 ;
        RECT 0.310 245.840 496.855 249.880 ;
        RECT 4.400 244.480 496.855 245.840 ;
        RECT 4.400 244.440 496.455 244.480 ;
        RECT 0.310 243.080 496.455 244.440 ;
        RECT 0.310 237.680 496.855 243.080 ;
        RECT 4.400 236.320 496.855 237.680 ;
        RECT 4.400 236.280 496.455 236.320 ;
        RECT 0.310 234.920 496.455 236.280 ;
        RECT 0.310 230.880 496.855 234.920 ;
        RECT 4.400 229.480 496.855 230.880 ;
        RECT 0.310 228.160 496.855 229.480 ;
        RECT 0.310 226.760 496.455 228.160 ;
        RECT 0.310 222.720 496.855 226.760 ;
        RECT 4.400 221.360 496.855 222.720 ;
        RECT 4.400 221.320 496.455 221.360 ;
        RECT 0.310 219.960 496.455 221.320 ;
        RECT 0.310 215.920 496.855 219.960 ;
        RECT 4.400 214.520 496.855 215.920 ;
        RECT 0.310 213.200 496.855 214.520 ;
        RECT 0.310 211.800 496.455 213.200 ;
        RECT 0.310 207.760 496.855 211.800 ;
        RECT 4.400 206.400 496.855 207.760 ;
        RECT 4.400 206.360 496.455 206.400 ;
        RECT 0.310 205.000 496.455 206.360 ;
        RECT 0.310 200.960 496.855 205.000 ;
        RECT 4.400 199.560 496.855 200.960 ;
        RECT 0.310 198.240 496.855 199.560 ;
        RECT 0.310 196.840 496.455 198.240 ;
        RECT 0.310 192.800 496.855 196.840 ;
        RECT 4.400 191.440 496.855 192.800 ;
        RECT 4.400 191.400 496.455 191.440 ;
        RECT 0.310 190.040 496.455 191.400 ;
        RECT 0.310 186.000 496.855 190.040 ;
        RECT 4.400 184.600 496.855 186.000 ;
        RECT 0.310 183.280 496.855 184.600 ;
        RECT 0.310 181.880 496.455 183.280 ;
        RECT 0.310 177.840 496.855 181.880 ;
        RECT 4.400 176.480 496.855 177.840 ;
        RECT 4.400 176.440 496.455 176.480 ;
        RECT 0.310 175.080 496.455 176.440 ;
        RECT 0.310 169.680 496.855 175.080 ;
        RECT 4.400 168.320 496.855 169.680 ;
        RECT 4.400 168.280 496.455 168.320 ;
        RECT 0.310 166.920 496.455 168.280 ;
        RECT 0.310 162.880 496.855 166.920 ;
        RECT 4.400 161.520 496.855 162.880 ;
        RECT 4.400 161.480 496.455 161.520 ;
        RECT 0.310 160.120 496.455 161.480 ;
        RECT 0.310 154.720 496.855 160.120 ;
        RECT 4.400 153.360 496.855 154.720 ;
        RECT 4.400 153.320 496.455 153.360 ;
        RECT 0.310 151.960 496.455 153.320 ;
        RECT 0.310 147.920 496.855 151.960 ;
        RECT 4.400 146.520 496.855 147.920 ;
        RECT 0.310 145.200 496.855 146.520 ;
        RECT 0.310 143.800 496.455 145.200 ;
        RECT 0.310 139.760 496.855 143.800 ;
        RECT 4.400 138.400 496.855 139.760 ;
        RECT 4.400 138.360 496.455 138.400 ;
        RECT 0.310 137.000 496.455 138.360 ;
        RECT 0.310 132.960 496.855 137.000 ;
        RECT 4.400 131.560 496.855 132.960 ;
        RECT 0.310 130.240 496.855 131.560 ;
        RECT 0.310 128.840 496.455 130.240 ;
        RECT 0.310 124.800 496.855 128.840 ;
        RECT 4.400 123.440 496.855 124.800 ;
        RECT 4.400 123.400 496.455 123.440 ;
        RECT 0.310 122.040 496.455 123.400 ;
        RECT 0.310 118.000 496.855 122.040 ;
        RECT 4.400 116.600 496.855 118.000 ;
        RECT 0.310 115.280 496.855 116.600 ;
        RECT 0.310 113.880 496.455 115.280 ;
        RECT 0.310 109.840 496.855 113.880 ;
        RECT 4.400 108.480 496.855 109.840 ;
        RECT 4.400 108.440 496.455 108.480 ;
        RECT 0.310 107.080 496.455 108.440 ;
        RECT 0.310 103.040 496.855 107.080 ;
        RECT 4.400 101.640 496.855 103.040 ;
        RECT 0.310 100.320 496.855 101.640 ;
        RECT 0.310 98.920 496.455 100.320 ;
        RECT 0.310 94.880 496.855 98.920 ;
        RECT 4.400 93.520 496.855 94.880 ;
        RECT 4.400 93.480 496.455 93.520 ;
        RECT 0.310 92.120 496.455 93.480 ;
        RECT 0.310 86.720 496.855 92.120 ;
        RECT 4.400 85.360 496.855 86.720 ;
        RECT 4.400 85.320 496.455 85.360 ;
        RECT 0.310 83.960 496.455 85.320 ;
        RECT 0.310 79.920 496.855 83.960 ;
        RECT 4.400 78.560 496.855 79.920 ;
        RECT 4.400 78.520 496.455 78.560 ;
        RECT 0.310 77.160 496.455 78.520 ;
        RECT 0.310 71.760 496.855 77.160 ;
        RECT 4.400 70.400 496.855 71.760 ;
        RECT 4.400 70.360 496.455 70.400 ;
        RECT 0.310 69.000 496.455 70.360 ;
        RECT 0.310 64.960 496.855 69.000 ;
        RECT 4.400 63.560 496.855 64.960 ;
        RECT 0.310 62.240 496.855 63.560 ;
        RECT 0.310 60.840 496.455 62.240 ;
        RECT 0.310 56.800 496.855 60.840 ;
        RECT 4.400 55.440 496.855 56.800 ;
        RECT 4.400 55.400 496.455 55.440 ;
        RECT 0.310 54.040 496.455 55.400 ;
        RECT 0.310 50.000 496.855 54.040 ;
        RECT 4.400 48.600 496.855 50.000 ;
        RECT 0.310 47.280 496.855 48.600 ;
        RECT 0.310 45.880 496.455 47.280 ;
        RECT 0.310 41.840 496.855 45.880 ;
        RECT 4.400 40.480 496.855 41.840 ;
        RECT 4.400 40.440 496.455 40.480 ;
        RECT 0.310 39.080 496.455 40.440 ;
        RECT 0.310 35.040 496.855 39.080 ;
        RECT 4.400 33.640 496.855 35.040 ;
        RECT 0.310 32.320 496.855 33.640 ;
        RECT 0.310 30.920 496.455 32.320 ;
        RECT 0.310 26.880 496.855 30.920 ;
        RECT 4.400 25.520 496.855 26.880 ;
        RECT 4.400 25.480 496.455 25.520 ;
        RECT 0.310 24.120 496.455 25.480 ;
        RECT 0.310 20.080 496.855 24.120 ;
        RECT 4.400 18.680 496.855 20.080 ;
        RECT 0.310 17.360 496.855 18.680 ;
        RECT 0.310 15.960 496.455 17.360 ;
        RECT 0.310 11.920 496.855 15.960 ;
        RECT 4.400 10.560 496.855 11.920 ;
        RECT 4.400 10.520 496.455 10.560 ;
        RECT 0.310 9.160 496.455 10.520 ;
        RECT 0.310 4.255 496.855 9.160 ;
      LAYER met4 ;
        RECT 15.935 10.640 483.440 500.720 ;
      LAYER met5 ;
        RECT 5.520 179.670 494.960 487.630 ;
  END
END mac_cluster
END LIBRARY

