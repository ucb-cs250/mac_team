`define MAC_SINGLE 0
`define MAC_DUAL 1
`define MAC_QUAD 2
