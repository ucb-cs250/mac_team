VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mac_cluster
  CLASS BLOCK ;
  FOREIGN mac_cluster ;
  ORIGIN 0.000 0.000 ;
  SIZE 505.140 BY 515.860 ;
  PIN A0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 188.690 511.860 188.970 515.860 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 274.760 505.140 275.360 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 425.130 511.860 425.410 515.860 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.330 511.860 204.610 515.860 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END A0[7]
  PIN A1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.570 511.860 178.850 515.860 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 473.320 505.140 473.920 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.970 511.860 266.250 515.860 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 290.810 511.860 291.090 515.860 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 511.860 18.770 515.860 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 276.090 511.860 276.370 515.860 ;
    END
  END A1[7]
  PIN A2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.490 511.860 455.770 515.860 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END A2[6]
  PIN A2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 450.200 505.140 450.800 ;
    END
  END A2[7]
  PIN A3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.210 511.860 240.490 515.860 ;
    END
  END A3[0]
  PIN A3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END A3[1]
  PIN A3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.130 511.860 471.410 515.860 ;
    END
  END A3[2]
  PIN A3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.930 511.860 209.210 515.860 ;
    END
  END A3[3]
  PIN A3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END A3[4]
  PIN A3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END A3[5]
  PIN A3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END A3[6]
  PIN A3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.010 511.860 70.290 515.860 ;
    END
  END A3[7]
  PIN B0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END B0[0]
  PIN B0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END B0[1]
  PIN B0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END B0[2]
  PIN B0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END B0[3]
  PIN B0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 221.720 505.140 222.320 ;
    END
  END B0[4]
  PIN B0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 229.170 511.860 229.450 515.860 ;
    END
  END B0[5]
  PIN B0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 511.860 75.810 515.860 ;
    END
  END B0[6]
  PIN B0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END B0[7]
  PIN B1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 147.290 511.860 147.570 515.860 ;
    END
  END B1[0]
  PIN B1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 374.040 505.140 374.640 ;
    END
  END B1[1]
  PIN B1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 153.720 505.140 154.320 ;
    END
  END B1[2]
  PIN B1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END B1[3]
  PIN B1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 378.210 511.860 378.490 515.860 ;
    END
  END B1[4]
  PIN B1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END B1[5]
  PIN B1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.410 511.860 157.690 515.860 ;
    END
  END B1[6]
  PIN B1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 244.840 505.140 245.440 ;
    END
  END B1[7]
  PIN B2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END B2[0]
  PIN B2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END B2[1]
  PIN B2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END B2[2]
  PIN B2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 115.640 505.140 116.240 ;
    END
  END B2[3]
  PIN B2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 162.930 511.860 163.210 515.860 ;
    END
  END B2[4]
  PIN B2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 511.860 24.290 515.860 ;
    END
  END B2[5]
  PIN B2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END B2[6]
  PIN B2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 282.920 505.140 283.520 ;
    END
  END B2[7]
  PIN B3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 77.560 505.140 78.160 ;
    END
  END B3[0]
  PIN B3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END B3[1]
  PIN B3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END B3[2]
  PIN B3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 488.280 505.140 488.880 ;
    END
  END B3[3]
  PIN B3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 214.920 505.140 215.520 ;
    END
  END B3[4]
  PIN B3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 511.860 29.810 515.860 ;
    END
  END B3[5]
  PIN B3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END B3[6]
  PIN B3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 107.480 505.140 108.080 ;
    END
  END B3[7]
  PIN cfg[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 260.450 511.860 260.730 515.860 ;
    END
  END cfg[0]
  PIN cfg[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END cfg[100]
  PIN cfg[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END cfg[101]
  PIN cfg[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END cfg[102]
  PIN cfg[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 511.860 50.050 515.860 ;
    END
  END cfg[103]
  PIN cfg[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END cfg[104]
  PIN cfg[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END cfg[105]
  PIN cfg[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 435.240 505.140 435.840 ;
    END
  END cfg[106]
  PIN cfg[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END cfg[107]
  PIN cfg[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END cfg[108]
  PIN cfg[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.410 511.860 111.690 515.860 ;
    END
  END cfg[109]
  PIN cfg[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END cfg[10]
  PIN cfg[110]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END cfg[110]
  PIN cfg[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END cfg[111]
  PIN cfg[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END cfg[112]
  PIN cfg[113]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 206.760 505.140 207.360 ;
    END
  END cfg[113]
  PIN cfg[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 253.000 505.140 253.600 ;
    END
  END cfg[114]
  PIN cfg[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.170 511.860 91.450 515.860 ;
    END
  END cfg[115]
  PIN cfg[116]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END cfg[116]
  PIN cfg[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 435.250 511.860 435.530 515.860 ;
    END
  END cfg[117]
  PIN cfg[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END cfg[118]
  PIN cfg[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END cfg[119]
  PIN cfg[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END cfg[11]
  PIN cfg[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.530 511.860 121.810 515.860 ;
    END
  END cfg[120]
  PIN cfg[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 24.520 505.140 25.120 ;
    END
  END cfg[121]
  PIN cfg[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END cfg[122]
  PIN cfg[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END cfg[123]
  PIN cfg[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 365.880 505.140 366.480 ;
    END
  END cfg[124]
  PIN cfg[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 511.860 34.410 515.860 ;
    END
  END cfg[125]
  PIN cfg[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 259.800 505.140 260.400 ;
    END
  END cfg[126]
  PIN cfg[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END cfg[127]
  PIN cfg[128]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END cfg[128]
  PIN cfg[129]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END cfg[129]
  PIN cfg[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END cfg[12]
  PIN cfg[130]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END cfg[130]
  PIN cfg[131]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.370 511.860 353.650 515.860 ;
    END
  END cfg[131]
  PIN cfg[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 327.610 511.860 327.890 515.860 ;
    END
  END cfg[13]
  PIN cfg[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END cfg[14]
  PIN cfg[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END cfg[15]
  PIN cfg[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END cfg[16]
  PIN cfg[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 296.330 511.860 296.610 515.860 ;
    END
  END cfg[17]
  PIN cfg[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 359.080 505.140 359.680 ;
    END
  END cfg[18]
  PIN cfg[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END cfg[19]
  PIN cfg[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END cfg[1]
  PIN cfg[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 214.450 511.860 214.730 515.860 ;
    END
  END cfg[20]
  PIN cfg[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 92.520 505.140 93.120 ;
    END
  END cfg[21]
  PIN cfg[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 176.840 505.140 177.440 ;
    END
  END cfg[22]
  PIN cfg[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END cfg[23]
  PIN cfg[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 16.360 505.140 16.960 ;
    END
  END cfg[24]
  PIN cfg[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END cfg[25]
  PIN cfg[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END cfg[26]
  PIN cfg[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 342.330 511.860 342.610 515.860 ;
    END
  END cfg[27]
  PIN cfg[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 439.850 511.860 440.130 515.860 ;
    END
  END cfg[28]
  PIN cfg[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END cfg[29]
  PIN cfg[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END cfg[2]
  PIN cfg[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END cfg[30]
  PIN cfg[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 321.000 505.140 321.600 ;
    END
  END cfg[31]
  PIN cfg[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 476.650 511.860 476.930 515.860 ;
    END
  END cfg[32]
  PIN cfg[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.930 511.860 255.210 515.860 ;
    END
  END cfg[33]
  PIN cfg[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END cfg[34]
  PIN cfg[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END cfg[35]
  PIN cfg[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END cfg[36]
  PIN cfg[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END cfg[37]
  PIN cfg[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 54.440 505.140 55.040 ;
    END
  END cfg[38]
  PIN cfg[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 389.000 505.140 389.600 ;
    END
  END cfg[39]
  PIN cfg[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 465.160 505.140 465.760 ;
    END
  END cfg[3]
  PIN cfg[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 480.330 0.000 480.610 4.000 ;
    END
  END cfg[40]
  PIN cfg[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 511.860 85.930 515.860 ;
    END
  END cfg[41]
  PIN cfg[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END cfg[42]
  PIN cfg[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END cfg[43]
  PIN cfg[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 130.600 505.140 131.200 ;
    END
  END cfg[44]
  PIN cfg[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END cfg[45]
  PIN cfg[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 412.120 505.140 412.720 ;
    END
  END cfg[46]
  PIN cfg[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.970 511.860 404.250 515.860 ;
    END
  END cfg[47]
  PIN cfg[48]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END cfg[48]
  PIN cfg[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 511.860 80.410 515.860 ;
    END
  END cfg[49]
  PIN cfg[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.050 511.860 173.330 515.860 ;
    END
  END cfg[4]
  PIN cfg[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END cfg[50]
  PIN cfg[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 465.610 511.860 465.890 515.860 ;
    END
  END cfg[51]
  PIN cfg[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END cfg[52]
  PIN cfg[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END cfg[53]
  PIN cfg[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END cfg[54]
  PIN cfg[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END cfg[55]
  PIN cfg[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END cfg[56]
  PIN cfg[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END cfg[57]
  PIN cfg[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.250 511.860 389.530 515.860 ;
    END
  END cfg[58]
  PIN cfg[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END cfg[59]
  PIN cfg[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 393.850 511.860 394.130 515.860 ;
    END
  END cfg[5]
  PIN cfg[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 495.080 505.140 495.680 ;
    END
  END cfg[60]
  PIN cfg[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 297.880 505.140 298.480 ;
    END
  END cfg[61]
  PIN cfg[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 301.850 511.860 302.130 515.860 ;
    END
  END cfg[62]
  PIN cfg[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 145.560 505.140 146.160 ;
    END
  END cfg[63]
  PIN cfg[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END cfg[64]
  PIN cfg[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END cfg[65]
  PIN cfg[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 511.860 106.170 515.860 ;
    END
  END cfg[66]
  PIN cfg[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 511.860 4.050 515.860 ;
    END
  END cfg[67]
  PIN cfg[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END cfg[68]
  PIN cfg[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END cfg[69]
  PIN cfg[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 306.450 511.860 306.730 515.860 ;
    END
  END cfg[6]
  PIN cfg[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END cfg[70]
  PIN cfg[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 161.880 505.140 162.480 ;
    END
  END cfg[71]
  PIN cfg[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END cfg[72]
  PIN cfg[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END cfg[73]
  PIN cfg[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 167.530 511.860 167.810 515.860 ;
    END
  END cfg[74]
  PIN cfg[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END cfg[75]
  PIN cfg[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END cfg[76]
  PIN cfg[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END cfg[77]
  PIN cfg[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 32.680 505.140 33.280 ;
    END
  END cfg[78]
  PIN cfg[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 409.490 511.860 409.770 515.860 ;
    END
  END cfg[79]
  PIN cfg[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END cfg[7]
  PIN cfg[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END cfg[80]
  PIN cfg[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END cfg[81]
  PIN cfg[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END cfg[82]
  PIN cfg[83]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END cfg[83]
  PIN cfg[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 510.040 505.140 510.640 ;
    END
  END cfg[84]
  PIN cfg[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 363.490 511.860 363.770 515.860 ;
    END
  END cfg[85]
  PIN cfg[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.090 511.860 322.370 515.860 ;
    END
  END cfg[86]
  PIN cfg[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 199.960 505.140 200.560 ;
    END
  END cfg[87]
  PIN cfg[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.730 511.860 338.010 515.860 ;
    END
  END cfg[88]
  PIN cfg[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END cfg[89]
  PIN cfg[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 335.960 505.140 336.560 ;
    END
  END cfg[8]
  PIN cfg[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END cfg[90]
  PIN cfg[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END cfg[91]
  PIN cfg[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END cfg[92]
  PIN cfg[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END cfg[93]
  PIN cfg[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END cfg[94]
  PIN cfg[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.930 511.860 117.210 515.860 ;
    END
  END cfg[95]
  PIN cfg[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 100.680 505.140 101.280 ;
    END
  END cfg[96]
  PIN cfg[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END cfg[97]
  PIN cfg[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END cfg[98]
  PIN cfg[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END cfg[99]
  PIN cfg[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 418.920 505.140 419.520 ;
    END
  END cfg[9]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 481.250 511.860 481.530 515.860 ;
    END
  END clk
  PIN cset
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 501.140 229.880 505.140 230.480 ;
    END
  END cset
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 280.690 511.860 280.970 515.860 ;
    END
  END en
  PIN out0[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END out0[0]
  PIN out0[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 419.610 511.860 419.890 515.860 ;
    END
  END out0[10]
  PIN out0[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 267.960 505.140 268.560 ;
    END
  END out0[11]
  PIN out0[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 427.080 505.140 427.680 ;
    END
  END out0[12]
  PIN out0[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 306.040 505.140 306.640 ;
    END
  END out0[13]
  PIN out0[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 123.800 505.140 124.400 ;
    END
  END out0[14]
  PIN out0[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.170 511.860 183.450 515.860 ;
    END
  END out0[15]
  PIN out0[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 142.690 511.860 142.970 515.860 ;
    END
  END out0[16]
  PIN out0[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.050 511.860 127.330 515.860 ;
    END
  END out0[17]
  PIN out0[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END out0[18]
  PIN out0[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END out0[19]
  PIN out0[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 344.120 505.140 344.720 ;
    END
  END out0[1]
  PIN out0[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END out0[20]
  PIN out0[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END out0[21]
  PIN out0[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END out0[22]
  PIN out0[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END out0[23]
  PIN out0[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 224.570 511.860 224.850 515.860 ;
    END
  END out0[24]
  PIN out0[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 383.730 511.860 384.010 515.860 ;
    END
  END out0[25]
  PIN out0[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 403.960 505.140 404.560 ;
    END
  END out0[26]
  PIN out0[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 457.000 505.140 457.600 ;
    END
  END out0[27]
  PIN out0[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 511.860 55.570 515.860 ;
    END
  END out0[28]
  PIN out0[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 327.800 505.140 328.400 ;
    END
  END out0[29]
  PIN out0[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 461.010 511.860 461.290 515.860 ;
    END
  END out0[2]
  PIN out0[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END out0[30]
  PIN out0[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END out0[31]
  PIN out0[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END out0[3]
  PIN out0[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 39.480 505.140 40.080 ;
    END
  END out0[4]
  PIN out0[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 382.200 505.140 382.800 ;
    END
  END out0[5]
  PIN out0[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.850 511.860 348.130 515.860 ;
    END
  END out0[6]
  PIN out0[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 312.840 505.140 313.440 ;
    END
  END out0[7]
  PIN out0[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END out0[8]
  PIN out0[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 491.370 511.860 491.650 515.860 ;
    END
  END out0[9]
  PIN out1[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 332.210 511.860 332.490 515.860 ;
    END
  END out1[0]
  PIN out1[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 350.920 505.140 351.520 ;
    END
  END out1[10]
  PIN out1[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 442.040 505.140 442.640 ;
    END
  END out1[11]
  PIN out1[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END out1[12]
  PIN out1[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END out1[13]
  PIN out1[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.250 511.860 44.530 515.860 ;
    END
  END out1[14]
  PIN out1[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 311.970 511.860 312.250 515.860 ;
    END
  END out1[15]
  PIN out1[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END out1[16]
  PIN out1[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 191.800 505.140 192.400 ;
    END
  END out1[17]
  PIN out1[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.650 511.860 39.930 515.860 ;
    END
  END out1[18]
  PIN out1[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END out1[19]
  PIN out1[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END out1[1]
  PIN out1[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 480.120 505.140 480.720 ;
    END
  END out1[20]
  PIN out1[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 429.730 511.860 430.010 515.860 ;
    END
  END out1[21]
  PIN out1[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END out1[22]
  PIN out1[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END out1[23]
  PIN out1[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.650 511.860 131.930 515.860 ;
    END
  END out1[24]
  PIN out1[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END out1[25]
  PIN out1[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END out1[26]
  PIN out1[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 486.770 511.860 487.050 515.860 ;
    END
  END out1[27]
  PIN out1[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 168.680 505.140 169.280 ;
    END
  END out1[28]
  PIN out1[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 4.000 ;
    END
  END out1[29]
  PIN out1[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END out1[2]
  PIN out1[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END out1[30]
  PIN out1[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 511.860 14.170 515.860 ;
    END
  END out1[31]
  PIN out1[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 70.760 505.140 71.360 ;
    END
  END out1[3]
  PIN out1[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END out1[4]
  PIN out1[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END out1[5]
  PIN out1[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END out1[6]
  PIN out1[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 183.640 505.140 184.240 ;
    END
  END out1[7]
  PIN out1[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 219.050 511.860 219.330 515.860 ;
    END
  END out1[8]
  PIN out1[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.170 511.860 137.450 515.860 ;
    END
  END out1[9]
  PIN out2[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END out2[0]
  PIN out2[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END out2[10]
  PIN out2[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 511.860 101.570 515.860 ;
    END
  END out2[11]
  PIN out2[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 138.760 505.140 139.360 ;
    END
  END out2[12]
  PIN out2[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END out2[13]
  PIN out2[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END out2[14]
  PIN out2[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 250.330 511.860 250.610 515.860 ;
    END
  END out2[15]
  PIN out2[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 316.570 511.860 316.850 515.860 ;
    END
  END out2[16]
  PIN out2[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END out2[17]
  PIN out2[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 397.160 505.140 397.760 ;
    END
  END out2[18]
  PIN out2[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END out2[19]
  PIN out2[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END out2[1]
  PIN out2[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 152.810 511.860 153.090 515.860 ;
    END
  END out2[20]
  PIN out2[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END out2[21]
  PIN out2[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 503.240 505.140 503.840 ;
    END
  END out2[22]
  PIN out2[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END out2[23]
  PIN out2[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 236.680 505.140 237.280 ;
    END
  END out2[24]
  PIN out2[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END out2[25]
  PIN out2[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 47.640 505.140 48.240 ;
    END
  END out2[26]
  PIN out2[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END out2[27]
  PIN out2[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 450.890 511.860 451.170 515.860 ;
    END
  END out2[28]
  PIN out2[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END out2[29]
  PIN out2[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 244.810 511.860 245.090 515.860 ;
    END
  END out2[2]
  PIN out2[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END out2[30]
  PIN out2[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END out2[31]
  PIN out2[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 511.860 65.690 515.860 ;
    END
  END out2[3]
  PIN out2[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 399.370 511.860 399.650 515.860 ;
    END
  END out2[4]
  PIN out2[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 193.290 511.860 193.570 515.860 ;
    END
  END out2[5]
  PIN out2[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END out2[6]
  PIN out2[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.810 511.860 199.090 515.860 ;
    END
  END out2[7]
  PIN out2[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END out2[8]
  PIN out2[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 62.600 505.140 63.200 ;
    END
  END out2[9]
  PIN out3[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END out3[0]
  PIN out3[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.370 511.860 445.650 515.860 ;
    END
  END out3[10]
  PIN out3[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 286.210 511.860 286.490 515.860 ;
    END
  END out3[11]
  PIN out3[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.970 511.860 358.250 515.860 ;
    END
  END out3[12]
  PIN out3[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END out3[13]
  PIN out3[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END out3[14]
  PIN out3[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 291.080 505.140 291.680 ;
    END
  END out3[15]
  PIN out3[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END out3[16]
  PIN out3[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END out3[17]
  PIN out3[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.090 511.860 368.370 515.860 ;
    END
  END out3[18]
  PIN out3[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 511.860 96.050 515.860 ;
    END
  END out3[19]
  PIN out3[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 511.860 60.170 515.860 ;
    END
  END out3[1]
  PIN out3[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END out3[20]
  PIN out3[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END out3[21]
  PIN out3[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END out3[22]
  PIN out3[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 270.570 511.860 270.850 515.860 ;
    END
  END out3[23]
  PIN out3[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END out3[24]
  PIN out3[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 85.720 505.140 86.320 ;
    END
  END out3[25]
  PIN out3[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END out3[26]
  PIN out3[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 511.860 8.650 515.860 ;
    END
  END out3[27]
  PIN out3[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 373.610 511.860 373.890 515.860 ;
    END
  END out3[28]
  PIN out3[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 415.010 511.860 415.290 515.860 ;
    END
  END out3[29]
  PIN out3[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END out3[2]
  PIN out3[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END out3[30]
  PIN out3[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END out3[31]
  PIN out3[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END out3[3]
  PIN out3[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END out3[4]
  PIN out3[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.690 511.860 234.970 515.860 ;
    END
  END out3[5]
  PIN out3[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END out3[6]
  PIN out3[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 501.140 9.560 505.140 10.160 ;
    END
  END out3[7]
  PIN out3[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END out3[8]
  PIN out3[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 496.890 511.860 497.170 515.860 ;
    END
  END out3[9]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END rst
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 499.560 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 499.560 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.065 10.795 499.560 503.285 ;
      LAYER met1 ;
        RECT 0.070 5.480 499.560 511.660 ;
      LAYER met2 ;
        RECT 0.100 511.580 3.490 511.860 ;
        RECT 4.330 511.580 8.090 511.860 ;
        RECT 8.930 511.580 13.610 511.860 ;
        RECT 14.450 511.580 18.210 511.860 ;
        RECT 19.050 511.580 23.730 511.860 ;
        RECT 24.570 511.580 29.250 511.860 ;
        RECT 30.090 511.580 33.850 511.860 ;
        RECT 34.690 511.580 39.370 511.860 ;
        RECT 40.210 511.580 43.970 511.860 ;
        RECT 44.810 511.580 49.490 511.860 ;
        RECT 50.330 511.580 55.010 511.860 ;
        RECT 55.850 511.580 59.610 511.860 ;
        RECT 60.450 511.580 65.130 511.860 ;
        RECT 65.970 511.580 69.730 511.860 ;
        RECT 70.570 511.580 75.250 511.860 ;
        RECT 76.090 511.580 79.850 511.860 ;
        RECT 80.690 511.580 85.370 511.860 ;
        RECT 86.210 511.580 90.890 511.860 ;
        RECT 91.730 511.580 95.490 511.860 ;
        RECT 96.330 511.580 101.010 511.860 ;
        RECT 101.850 511.580 105.610 511.860 ;
        RECT 106.450 511.580 111.130 511.860 ;
        RECT 111.970 511.580 116.650 511.860 ;
        RECT 117.490 511.580 121.250 511.860 ;
        RECT 122.090 511.580 126.770 511.860 ;
        RECT 127.610 511.580 131.370 511.860 ;
        RECT 132.210 511.580 136.890 511.860 ;
        RECT 137.730 511.580 142.410 511.860 ;
        RECT 143.250 511.580 147.010 511.860 ;
        RECT 147.850 511.580 152.530 511.860 ;
        RECT 153.370 511.580 157.130 511.860 ;
        RECT 157.970 511.580 162.650 511.860 ;
        RECT 163.490 511.580 167.250 511.860 ;
        RECT 168.090 511.580 172.770 511.860 ;
        RECT 173.610 511.580 178.290 511.860 ;
        RECT 179.130 511.580 182.890 511.860 ;
        RECT 183.730 511.580 188.410 511.860 ;
        RECT 189.250 511.580 193.010 511.860 ;
        RECT 193.850 511.580 198.530 511.860 ;
        RECT 199.370 511.580 204.050 511.860 ;
        RECT 204.890 511.580 208.650 511.860 ;
        RECT 209.490 511.580 214.170 511.860 ;
        RECT 215.010 511.580 218.770 511.860 ;
        RECT 219.610 511.580 224.290 511.860 ;
        RECT 225.130 511.580 228.890 511.860 ;
        RECT 229.730 511.580 234.410 511.860 ;
        RECT 235.250 511.580 239.930 511.860 ;
        RECT 240.770 511.580 244.530 511.860 ;
        RECT 245.370 511.580 250.050 511.860 ;
        RECT 250.890 511.580 254.650 511.860 ;
        RECT 255.490 511.580 260.170 511.860 ;
        RECT 261.010 511.580 265.690 511.860 ;
        RECT 266.530 511.580 270.290 511.860 ;
        RECT 271.130 511.580 275.810 511.860 ;
        RECT 276.650 511.580 280.410 511.860 ;
        RECT 281.250 511.580 285.930 511.860 ;
        RECT 286.770 511.580 290.530 511.860 ;
        RECT 291.370 511.580 296.050 511.860 ;
        RECT 296.890 511.580 301.570 511.860 ;
        RECT 302.410 511.580 306.170 511.860 ;
        RECT 307.010 511.580 311.690 511.860 ;
        RECT 312.530 511.580 316.290 511.860 ;
        RECT 317.130 511.580 321.810 511.860 ;
        RECT 322.650 511.580 327.330 511.860 ;
        RECT 328.170 511.580 331.930 511.860 ;
        RECT 332.770 511.580 337.450 511.860 ;
        RECT 338.290 511.580 342.050 511.860 ;
        RECT 342.890 511.580 347.570 511.860 ;
        RECT 348.410 511.580 353.090 511.860 ;
        RECT 353.930 511.580 357.690 511.860 ;
        RECT 358.530 511.580 363.210 511.860 ;
        RECT 364.050 511.580 367.810 511.860 ;
        RECT 368.650 511.580 373.330 511.860 ;
        RECT 374.170 511.580 377.930 511.860 ;
        RECT 378.770 511.580 383.450 511.860 ;
        RECT 384.290 511.580 388.970 511.860 ;
        RECT 389.810 511.580 393.570 511.860 ;
        RECT 394.410 511.580 399.090 511.860 ;
        RECT 399.930 511.580 403.690 511.860 ;
        RECT 404.530 511.580 409.210 511.860 ;
        RECT 410.050 511.580 414.730 511.860 ;
        RECT 415.570 511.580 419.330 511.860 ;
        RECT 420.170 511.580 424.850 511.860 ;
        RECT 425.690 511.580 429.450 511.860 ;
        RECT 430.290 511.580 434.970 511.860 ;
        RECT 435.810 511.580 439.570 511.860 ;
        RECT 440.410 511.580 445.090 511.860 ;
        RECT 445.930 511.580 450.610 511.860 ;
        RECT 451.450 511.580 455.210 511.860 ;
        RECT 456.050 511.580 460.730 511.860 ;
        RECT 461.570 511.580 465.330 511.860 ;
        RECT 466.170 511.580 470.850 511.860 ;
        RECT 471.690 511.580 476.370 511.860 ;
        RECT 477.210 511.580 480.970 511.860 ;
        RECT 481.810 511.580 486.490 511.860 ;
        RECT 487.330 511.580 491.090 511.860 ;
        RECT 491.930 511.580 496.610 511.860 ;
        RECT 497.450 511.580 500.780 511.860 ;
        RECT 0.100 4.280 500.780 511.580 ;
        RECT 0.100 4.000 2.570 4.280 ;
        RECT 3.410 4.000 7.170 4.280 ;
        RECT 8.010 4.000 12.690 4.280 ;
        RECT 13.530 4.000 17.290 4.280 ;
        RECT 18.130 4.000 22.810 4.280 ;
        RECT 23.650 4.000 27.410 4.280 ;
        RECT 28.250 4.000 32.930 4.280 ;
        RECT 33.770 4.000 38.450 4.280 ;
        RECT 39.290 4.000 43.050 4.280 ;
        RECT 43.890 4.000 48.570 4.280 ;
        RECT 49.410 4.000 53.170 4.280 ;
        RECT 54.010 4.000 58.690 4.280 ;
        RECT 59.530 4.000 64.210 4.280 ;
        RECT 65.050 4.000 68.810 4.280 ;
        RECT 69.650 4.000 74.330 4.280 ;
        RECT 75.170 4.000 78.930 4.280 ;
        RECT 79.770 4.000 84.450 4.280 ;
        RECT 85.290 4.000 89.050 4.280 ;
        RECT 89.890 4.000 94.570 4.280 ;
        RECT 95.410 4.000 100.090 4.280 ;
        RECT 100.930 4.000 104.690 4.280 ;
        RECT 105.530 4.000 110.210 4.280 ;
        RECT 111.050 4.000 114.810 4.280 ;
        RECT 115.650 4.000 120.330 4.280 ;
        RECT 121.170 4.000 125.850 4.280 ;
        RECT 126.690 4.000 130.450 4.280 ;
        RECT 131.290 4.000 135.970 4.280 ;
        RECT 136.810 4.000 140.570 4.280 ;
        RECT 141.410 4.000 146.090 4.280 ;
        RECT 146.930 4.000 150.690 4.280 ;
        RECT 151.530 4.000 156.210 4.280 ;
        RECT 157.050 4.000 161.730 4.280 ;
        RECT 162.570 4.000 166.330 4.280 ;
        RECT 167.170 4.000 171.850 4.280 ;
        RECT 172.690 4.000 176.450 4.280 ;
        RECT 177.290 4.000 181.970 4.280 ;
        RECT 182.810 4.000 187.490 4.280 ;
        RECT 188.330 4.000 192.090 4.280 ;
        RECT 192.930 4.000 197.610 4.280 ;
        RECT 198.450 4.000 202.210 4.280 ;
        RECT 203.050 4.000 207.730 4.280 ;
        RECT 208.570 4.000 212.330 4.280 ;
        RECT 213.170 4.000 217.850 4.280 ;
        RECT 218.690 4.000 223.370 4.280 ;
        RECT 224.210 4.000 227.970 4.280 ;
        RECT 228.810 4.000 233.490 4.280 ;
        RECT 234.330 4.000 238.090 4.280 ;
        RECT 238.930 4.000 243.610 4.280 ;
        RECT 244.450 4.000 249.130 4.280 ;
        RECT 249.970 4.000 253.730 4.280 ;
        RECT 254.570 4.000 259.250 4.280 ;
        RECT 260.090 4.000 263.850 4.280 ;
        RECT 264.690 4.000 269.370 4.280 ;
        RECT 270.210 4.000 274.890 4.280 ;
        RECT 275.730 4.000 279.490 4.280 ;
        RECT 280.330 4.000 285.010 4.280 ;
        RECT 285.850 4.000 289.610 4.280 ;
        RECT 290.450 4.000 295.130 4.280 ;
        RECT 295.970 4.000 299.730 4.280 ;
        RECT 300.570 4.000 305.250 4.280 ;
        RECT 306.090 4.000 310.770 4.280 ;
        RECT 311.610 4.000 315.370 4.280 ;
        RECT 316.210 4.000 320.890 4.280 ;
        RECT 321.730 4.000 325.490 4.280 ;
        RECT 326.330 4.000 331.010 4.280 ;
        RECT 331.850 4.000 336.530 4.280 ;
        RECT 337.370 4.000 341.130 4.280 ;
        RECT 341.970 4.000 346.650 4.280 ;
        RECT 347.490 4.000 351.250 4.280 ;
        RECT 352.090 4.000 356.770 4.280 ;
        RECT 357.610 4.000 361.370 4.280 ;
        RECT 362.210 4.000 366.890 4.280 ;
        RECT 367.730 4.000 372.410 4.280 ;
        RECT 373.250 4.000 377.010 4.280 ;
        RECT 377.850 4.000 382.530 4.280 ;
        RECT 383.370 4.000 387.130 4.280 ;
        RECT 387.970 4.000 392.650 4.280 ;
        RECT 393.490 4.000 398.170 4.280 ;
        RECT 399.010 4.000 402.770 4.280 ;
        RECT 403.610 4.000 408.290 4.280 ;
        RECT 409.130 4.000 412.890 4.280 ;
        RECT 413.730 4.000 418.410 4.280 ;
        RECT 419.250 4.000 423.010 4.280 ;
        RECT 423.850 4.000 428.530 4.280 ;
        RECT 429.370 4.000 434.050 4.280 ;
        RECT 434.890 4.000 438.650 4.280 ;
        RECT 439.490 4.000 444.170 4.280 ;
        RECT 445.010 4.000 448.770 4.280 ;
        RECT 449.610 4.000 454.290 4.280 ;
        RECT 455.130 4.000 459.810 4.280 ;
        RECT 460.650 4.000 464.410 4.280 ;
        RECT 465.250 4.000 469.930 4.280 ;
        RECT 470.770 4.000 474.530 4.280 ;
        RECT 475.370 4.000 480.050 4.280 ;
        RECT 480.890 4.000 485.570 4.280 ;
        RECT 486.410 4.000 490.170 4.280 ;
        RECT 491.010 4.000 495.690 4.280 ;
        RECT 496.530 4.000 500.290 4.280 ;
      LAYER met3 ;
        RECT 4.000 509.640 500.740 510.505 ;
        RECT 4.000 505.600 501.140 509.640 ;
        RECT 4.400 504.240 501.140 505.600 ;
        RECT 4.400 504.200 500.740 504.240 ;
        RECT 4.000 502.840 500.740 504.200 ;
        RECT 4.000 498.800 501.140 502.840 ;
        RECT 4.400 497.400 501.140 498.800 ;
        RECT 4.000 496.080 501.140 497.400 ;
        RECT 4.000 494.680 500.740 496.080 ;
        RECT 4.000 490.640 501.140 494.680 ;
        RECT 4.400 489.280 501.140 490.640 ;
        RECT 4.400 489.240 500.740 489.280 ;
        RECT 4.000 487.880 500.740 489.240 ;
        RECT 4.000 482.480 501.140 487.880 ;
        RECT 4.400 481.120 501.140 482.480 ;
        RECT 4.400 481.080 500.740 481.120 ;
        RECT 4.000 479.720 500.740 481.080 ;
        RECT 4.000 475.680 501.140 479.720 ;
        RECT 4.400 474.320 501.140 475.680 ;
        RECT 4.400 474.280 500.740 474.320 ;
        RECT 4.000 472.920 500.740 474.280 ;
        RECT 4.000 467.520 501.140 472.920 ;
        RECT 4.400 466.160 501.140 467.520 ;
        RECT 4.400 466.120 500.740 466.160 ;
        RECT 4.000 464.760 500.740 466.120 ;
        RECT 4.000 460.720 501.140 464.760 ;
        RECT 4.400 459.320 501.140 460.720 ;
        RECT 4.000 458.000 501.140 459.320 ;
        RECT 4.000 456.600 500.740 458.000 ;
        RECT 4.000 452.560 501.140 456.600 ;
        RECT 4.400 451.200 501.140 452.560 ;
        RECT 4.400 451.160 500.740 451.200 ;
        RECT 4.000 449.800 500.740 451.160 ;
        RECT 4.000 444.400 501.140 449.800 ;
        RECT 4.400 443.040 501.140 444.400 ;
        RECT 4.400 443.000 500.740 443.040 ;
        RECT 4.000 441.640 500.740 443.000 ;
        RECT 4.000 437.600 501.140 441.640 ;
        RECT 4.400 436.240 501.140 437.600 ;
        RECT 4.400 436.200 500.740 436.240 ;
        RECT 4.000 434.840 500.740 436.200 ;
        RECT 4.000 429.440 501.140 434.840 ;
        RECT 4.400 428.080 501.140 429.440 ;
        RECT 4.400 428.040 500.740 428.080 ;
        RECT 4.000 426.680 500.740 428.040 ;
        RECT 4.000 422.640 501.140 426.680 ;
        RECT 4.400 421.240 501.140 422.640 ;
        RECT 4.000 419.920 501.140 421.240 ;
        RECT 4.000 418.520 500.740 419.920 ;
        RECT 4.000 414.480 501.140 418.520 ;
        RECT 4.400 413.120 501.140 414.480 ;
        RECT 4.400 413.080 500.740 413.120 ;
        RECT 4.000 411.720 500.740 413.080 ;
        RECT 4.000 407.680 501.140 411.720 ;
        RECT 4.400 406.280 501.140 407.680 ;
        RECT 4.000 404.960 501.140 406.280 ;
        RECT 4.000 403.560 500.740 404.960 ;
        RECT 4.000 399.520 501.140 403.560 ;
        RECT 4.400 398.160 501.140 399.520 ;
        RECT 4.400 398.120 500.740 398.160 ;
        RECT 4.000 396.760 500.740 398.120 ;
        RECT 4.000 391.360 501.140 396.760 ;
        RECT 4.400 390.000 501.140 391.360 ;
        RECT 4.400 389.960 500.740 390.000 ;
        RECT 4.000 388.600 500.740 389.960 ;
        RECT 4.000 384.560 501.140 388.600 ;
        RECT 4.400 383.200 501.140 384.560 ;
        RECT 4.400 383.160 500.740 383.200 ;
        RECT 4.000 381.800 500.740 383.160 ;
        RECT 4.000 376.400 501.140 381.800 ;
        RECT 4.400 375.040 501.140 376.400 ;
        RECT 4.400 375.000 500.740 375.040 ;
        RECT 4.000 373.640 500.740 375.000 ;
        RECT 4.000 369.600 501.140 373.640 ;
        RECT 4.400 368.200 501.140 369.600 ;
        RECT 4.000 366.880 501.140 368.200 ;
        RECT 4.000 365.480 500.740 366.880 ;
        RECT 4.000 361.440 501.140 365.480 ;
        RECT 4.400 360.080 501.140 361.440 ;
        RECT 4.400 360.040 500.740 360.080 ;
        RECT 4.000 358.680 500.740 360.040 ;
        RECT 4.000 353.280 501.140 358.680 ;
        RECT 4.400 351.920 501.140 353.280 ;
        RECT 4.400 351.880 500.740 351.920 ;
        RECT 4.000 350.520 500.740 351.880 ;
        RECT 4.000 346.480 501.140 350.520 ;
        RECT 4.400 345.120 501.140 346.480 ;
        RECT 4.400 345.080 500.740 345.120 ;
        RECT 4.000 343.720 500.740 345.080 ;
        RECT 4.000 338.320 501.140 343.720 ;
        RECT 4.400 336.960 501.140 338.320 ;
        RECT 4.400 336.920 500.740 336.960 ;
        RECT 4.000 335.560 500.740 336.920 ;
        RECT 4.000 331.520 501.140 335.560 ;
        RECT 4.400 330.120 501.140 331.520 ;
        RECT 4.000 328.800 501.140 330.120 ;
        RECT 4.000 327.400 500.740 328.800 ;
        RECT 4.000 323.360 501.140 327.400 ;
        RECT 4.400 322.000 501.140 323.360 ;
        RECT 4.400 321.960 500.740 322.000 ;
        RECT 4.000 320.600 500.740 321.960 ;
        RECT 4.000 315.200 501.140 320.600 ;
        RECT 4.400 313.840 501.140 315.200 ;
        RECT 4.400 313.800 500.740 313.840 ;
        RECT 4.000 312.440 500.740 313.800 ;
        RECT 4.000 308.400 501.140 312.440 ;
        RECT 4.400 307.040 501.140 308.400 ;
        RECT 4.400 307.000 500.740 307.040 ;
        RECT 4.000 305.640 500.740 307.000 ;
        RECT 4.000 300.240 501.140 305.640 ;
        RECT 4.400 298.880 501.140 300.240 ;
        RECT 4.400 298.840 500.740 298.880 ;
        RECT 4.000 297.480 500.740 298.840 ;
        RECT 4.000 293.440 501.140 297.480 ;
        RECT 4.400 292.080 501.140 293.440 ;
        RECT 4.400 292.040 500.740 292.080 ;
        RECT 4.000 290.680 500.740 292.040 ;
        RECT 4.000 285.280 501.140 290.680 ;
        RECT 4.400 283.920 501.140 285.280 ;
        RECT 4.400 283.880 500.740 283.920 ;
        RECT 4.000 282.520 500.740 283.880 ;
        RECT 4.000 278.480 501.140 282.520 ;
        RECT 4.400 277.080 501.140 278.480 ;
        RECT 4.000 275.760 501.140 277.080 ;
        RECT 4.000 274.360 500.740 275.760 ;
        RECT 4.000 270.320 501.140 274.360 ;
        RECT 4.400 268.960 501.140 270.320 ;
        RECT 4.400 268.920 500.740 268.960 ;
        RECT 4.000 267.560 500.740 268.920 ;
        RECT 4.000 262.160 501.140 267.560 ;
        RECT 4.400 260.800 501.140 262.160 ;
        RECT 4.400 260.760 500.740 260.800 ;
        RECT 4.000 259.400 500.740 260.760 ;
        RECT 4.000 255.360 501.140 259.400 ;
        RECT 4.400 254.000 501.140 255.360 ;
        RECT 4.400 253.960 500.740 254.000 ;
        RECT 4.000 252.600 500.740 253.960 ;
        RECT 4.000 247.200 501.140 252.600 ;
        RECT 4.400 245.840 501.140 247.200 ;
        RECT 4.400 245.800 500.740 245.840 ;
        RECT 4.000 244.440 500.740 245.800 ;
        RECT 4.000 240.400 501.140 244.440 ;
        RECT 4.400 239.000 501.140 240.400 ;
        RECT 4.000 237.680 501.140 239.000 ;
        RECT 4.000 236.280 500.740 237.680 ;
        RECT 4.000 232.240 501.140 236.280 ;
        RECT 4.400 230.880 501.140 232.240 ;
        RECT 4.400 230.840 500.740 230.880 ;
        RECT 4.000 229.480 500.740 230.840 ;
        RECT 4.000 224.080 501.140 229.480 ;
        RECT 4.400 222.720 501.140 224.080 ;
        RECT 4.400 222.680 500.740 222.720 ;
        RECT 4.000 221.320 500.740 222.680 ;
        RECT 4.000 217.280 501.140 221.320 ;
        RECT 4.400 215.920 501.140 217.280 ;
        RECT 4.400 215.880 500.740 215.920 ;
        RECT 4.000 214.520 500.740 215.880 ;
        RECT 4.000 209.120 501.140 214.520 ;
        RECT 4.400 207.760 501.140 209.120 ;
        RECT 4.400 207.720 500.740 207.760 ;
        RECT 4.000 206.360 500.740 207.720 ;
        RECT 4.000 202.320 501.140 206.360 ;
        RECT 4.400 200.960 501.140 202.320 ;
        RECT 4.400 200.920 500.740 200.960 ;
        RECT 4.000 199.560 500.740 200.920 ;
        RECT 4.000 194.160 501.140 199.560 ;
        RECT 4.400 192.800 501.140 194.160 ;
        RECT 4.400 192.760 500.740 192.800 ;
        RECT 4.000 191.400 500.740 192.760 ;
        RECT 4.000 187.360 501.140 191.400 ;
        RECT 4.400 185.960 501.140 187.360 ;
        RECT 4.000 184.640 501.140 185.960 ;
        RECT 4.000 183.240 500.740 184.640 ;
        RECT 4.000 179.200 501.140 183.240 ;
        RECT 4.400 177.840 501.140 179.200 ;
        RECT 4.400 177.800 500.740 177.840 ;
        RECT 4.000 176.440 500.740 177.800 ;
        RECT 4.000 171.040 501.140 176.440 ;
        RECT 4.400 169.680 501.140 171.040 ;
        RECT 4.400 169.640 500.740 169.680 ;
        RECT 4.000 168.280 500.740 169.640 ;
        RECT 4.000 164.240 501.140 168.280 ;
        RECT 4.400 162.880 501.140 164.240 ;
        RECT 4.400 162.840 500.740 162.880 ;
        RECT 4.000 161.480 500.740 162.840 ;
        RECT 4.000 156.080 501.140 161.480 ;
        RECT 4.400 154.720 501.140 156.080 ;
        RECT 4.400 154.680 500.740 154.720 ;
        RECT 4.000 153.320 500.740 154.680 ;
        RECT 4.000 149.280 501.140 153.320 ;
        RECT 4.400 147.880 501.140 149.280 ;
        RECT 4.000 146.560 501.140 147.880 ;
        RECT 4.000 145.160 500.740 146.560 ;
        RECT 4.000 141.120 501.140 145.160 ;
        RECT 4.400 139.760 501.140 141.120 ;
        RECT 4.400 139.720 500.740 139.760 ;
        RECT 4.000 138.360 500.740 139.720 ;
        RECT 4.000 132.960 501.140 138.360 ;
        RECT 4.400 131.600 501.140 132.960 ;
        RECT 4.400 131.560 500.740 131.600 ;
        RECT 4.000 130.200 500.740 131.560 ;
        RECT 4.000 126.160 501.140 130.200 ;
        RECT 4.400 124.800 501.140 126.160 ;
        RECT 4.400 124.760 500.740 124.800 ;
        RECT 4.000 123.400 500.740 124.760 ;
        RECT 4.000 118.000 501.140 123.400 ;
        RECT 4.400 116.640 501.140 118.000 ;
        RECT 4.400 116.600 500.740 116.640 ;
        RECT 4.000 115.240 500.740 116.600 ;
        RECT 4.000 111.200 501.140 115.240 ;
        RECT 4.400 109.800 501.140 111.200 ;
        RECT 4.000 108.480 501.140 109.800 ;
        RECT 4.000 107.080 500.740 108.480 ;
        RECT 4.000 103.040 501.140 107.080 ;
        RECT 4.400 101.680 501.140 103.040 ;
        RECT 4.400 101.640 500.740 101.680 ;
        RECT 4.000 100.280 500.740 101.640 ;
        RECT 4.000 96.240 501.140 100.280 ;
        RECT 4.400 94.840 501.140 96.240 ;
        RECT 4.000 93.520 501.140 94.840 ;
        RECT 4.000 92.120 500.740 93.520 ;
        RECT 4.000 88.080 501.140 92.120 ;
        RECT 4.400 86.720 501.140 88.080 ;
        RECT 4.400 86.680 500.740 86.720 ;
        RECT 4.000 85.320 500.740 86.680 ;
        RECT 4.000 79.920 501.140 85.320 ;
        RECT 4.400 78.560 501.140 79.920 ;
        RECT 4.400 78.520 500.740 78.560 ;
        RECT 4.000 77.160 500.740 78.520 ;
        RECT 4.000 73.120 501.140 77.160 ;
        RECT 4.400 71.760 501.140 73.120 ;
        RECT 4.400 71.720 500.740 71.760 ;
        RECT 4.000 70.360 500.740 71.720 ;
        RECT 4.000 64.960 501.140 70.360 ;
        RECT 4.400 63.600 501.140 64.960 ;
        RECT 4.400 63.560 500.740 63.600 ;
        RECT 4.000 62.200 500.740 63.560 ;
        RECT 4.000 58.160 501.140 62.200 ;
        RECT 4.400 56.760 501.140 58.160 ;
        RECT 4.000 55.440 501.140 56.760 ;
        RECT 4.000 54.040 500.740 55.440 ;
        RECT 4.000 50.000 501.140 54.040 ;
        RECT 4.400 48.640 501.140 50.000 ;
        RECT 4.400 48.600 500.740 48.640 ;
        RECT 4.000 47.240 500.740 48.600 ;
        RECT 4.000 41.840 501.140 47.240 ;
        RECT 4.400 40.480 501.140 41.840 ;
        RECT 4.400 40.440 500.740 40.480 ;
        RECT 4.000 39.080 500.740 40.440 ;
        RECT 4.000 35.040 501.140 39.080 ;
        RECT 4.400 33.680 501.140 35.040 ;
        RECT 4.400 33.640 500.740 33.680 ;
        RECT 4.000 32.280 500.740 33.640 ;
        RECT 4.000 26.880 501.140 32.280 ;
        RECT 4.400 25.520 501.140 26.880 ;
        RECT 4.400 25.480 500.740 25.520 ;
        RECT 4.000 24.120 500.740 25.480 ;
        RECT 4.000 20.080 501.140 24.120 ;
        RECT 4.400 18.680 501.140 20.080 ;
        RECT 4.000 17.360 501.140 18.680 ;
        RECT 4.000 15.960 500.740 17.360 ;
        RECT 4.000 11.920 501.140 15.960 ;
        RECT 4.400 10.560 501.140 11.920 ;
        RECT 4.400 10.520 500.740 10.560 ;
        RECT 4.000 9.160 500.740 10.520 ;
        RECT 4.000 4.255 501.140 9.160 ;
      LAYER met4 ;
        RECT 19.615 10.640 486.385 503.705 ;
      LAYER met5 ;
        RECT 5.520 179.670 499.560 487.630 ;
  END
END mac_cluster
END LIBRARY

