VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mac_cluster
  CLASS BLOCK ;
  FOREIGN mac_cluster ;
  ORIGIN 0.000 0.000 ;
  SIZE 479.755 BY 490.475 ;
  PIN A0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.490 486.475 179.770 490.475 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 262.520 479.755 263.120 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.970 486.475 404.250 490.475 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.290 486.475 193.570 490.475 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END A0[7]
  PIN A1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.370 486.475 169.650 490.475 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 450.200 479.755 450.800 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 252.170 486.475 252.450 490.475 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 277.010 486.475 277.290 490.475 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 486.475 17.850 490.475 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 262.290 486.475 262.570 490.475 ;
    END
  END A1[7]
  PIN A2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 433.410 486.475 433.690 490.475 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END A2[6]
  PIN A2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 428.440 479.755 429.040 ;
    END
  END A2[7]
  PIN A3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.250 486.475 228.530 490.475 ;
    END
  END A3[0]
  PIN A3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END A3[1]
  PIN A3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 448.130 486.475 448.410 490.475 ;
    END
  END A3[2]
  PIN A3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 198.810 486.475 199.090 490.475 ;
    END
  END A3[3]
  PIN A3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END A3[4]
  PIN A3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END A3[5]
  PIN A3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END A3[6]
  PIN A3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.330 486.475 66.610 490.475 ;
    END
  END A3[7]
  PIN B0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END B0[0]
  PIN B0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END B0[1]
  PIN B0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END B0[2]
  PIN B0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END B0[3]
  PIN B0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 212.200 479.755 212.800 ;
    END
  END B0[4]
  PIN B0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.130 486.475 218.410 490.475 ;
    END
  END B0[5]
  PIN B0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 486.475 72.130 490.475 ;
    END
  END B0[6]
  PIN B0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END B0[7]
  PIN B1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.930 486.475 140.210 490.475 ;
    END
  END B1[0]
  PIN B1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 356.360 479.755 356.960 ;
    END
  END B1[1]
  PIN B1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 146.920 479.755 147.520 ;
    END
  END B1[2]
  PIN B1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END B1[3]
  PIN B1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 359.810 486.475 360.090 490.475 ;
    END
  END B1[4]
  PIN B1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END B1[5]
  PIN B1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.050 486.475 150.330 490.475 ;
    END
  END B1[6]
  PIN B1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 233.960 479.755 234.560 ;
    END
  END B1[7]
  PIN B2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END B2[0]
  PIN B2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END B2[1]
  PIN B2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END B2[2]
  PIN B2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 110.200 479.755 110.800 ;
    END
  END B2[3]
  PIN B2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.650 486.475 154.930 490.475 ;
    END
  END B2[4]
  PIN B2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 486.475 23.370 490.475 ;
    END
  END B2[5]
  PIN B2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END B2[6]
  PIN B2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 269.320 479.755 269.920 ;
    END
  END B2[7]
  PIN B3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 74.840 479.755 75.440 ;
    END
  END B3[0]
  PIN B3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END B3[1]
  PIN B3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END B3[2]
  PIN B3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 465.160 479.755 465.760 ;
    END
  END B3[3]
  PIN B3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 204.040 479.755 204.640 ;
    END
  END B3[4]
  PIN B3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.690 486.475 27.970 490.475 ;
    END
  END B3[5]
  PIN B3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END B3[6]
  PIN B3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 103.400 479.755 104.000 ;
    END
  END B3[7]
  PIN cfg[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.570 486.475 247.850 490.475 ;
    END
  END cfg[0]
  PIN cfg[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END cfg[100]
  PIN cfg[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END cfg[101]
  PIN cfg[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END cfg[102]
  PIN cfg[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 486.475 47.290 490.475 ;
    END
  END cfg[103]
  PIN cfg[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END cfg[104]
  PIN cfg[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END cfg[105]
  PIN cfg[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 413.480 479.755 414.080 ;
    END
  END cfg[106]
  PIN cfg[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END cfg[107]
  PIN cfg[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END cfg[108]
  PIN cfg[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 486.475 106.170 490.475 ;
    END
  END cfg[109]
  PIN cfg[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END cfg[10]
  PIN cfg[110]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END cfg[110]
  PIN cfg[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END cfg[111]
  PIN cfg[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END cfg[112]
  PIN cfg[113]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 197.240 479.755 197.840 ;
    END
  END cfg[113]
  PIN cfg[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 240.760 479.755 241.360 ;
    END
  END cfg[114]
  PIN cfg[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.570 486.475 86.850 490.475 ;
    END
  END cfg[115]
  PIN cfg[116]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END cfg[116]
  PIN cfg[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 413.170 486.475 413.450 490.475 ;
    END
  END cfg[117]
  PIN cfg[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END cfg[118]
  PIN cfg[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END cfg[119]
  PIN cfg[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END cfg[11]
  PIN cfg[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 486.475 115.370 490.475 ;
    END
  END cfg[120]
  PIN cfg[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 24.520 479.755 25.120 ;
    END
  END cfg[121]
  PIN cfg[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END cfg[122]
  PIN cfg[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END cfg[123]
  PIN cfg[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 349.560 479.755 350.160 ;
    END
  END cfg[124]
  PIN cfg[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 486.475 32.570 490.475 ;
    END
  END cfg[125]
  PIN cfg[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 247.560 479.755 248.160 ;
    END
  END cfg[126]
  PIN cfg[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END cfg[127]
  PIN cfg[128]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END cfg[128]
  PIN cfg[129]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END cfg[129]
  PIN cfg[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END cfg[12]
  PIN cfg[130]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END cfg[130]
  PIN cfg[131]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.970 486.475 335.250 490.475 ;
    END
  END cfg[131]
  PIN cfg[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.050 486.475 311.330 490.475 ;
    END
  END cfg[13]
  PIN cfg[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END cfg[14]
  PIN cfg[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END cfg[15]
  PIN cfg[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END cfg[16]
  PIN cfg[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.610 486.475 281.890 490.475 ;
    END
  END cfg[17]
  PIN cfg[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 341.400 479.755 342.000 ;
    END
  END cfg[18]
  PIN cfg[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END cfg[19]
  PIN cfg[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END cfg[1]
  PIN cfg[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 203.410 486.475 203.690 490.475 ;
    END
  END cfg[20]
  PIN cfg[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 88.440 479.755 89.040 ;
    END
  END cfg[21]
  PIN cfg[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 168.680 479.755 169.280 ;
    END
  END cfg[22]
  PIN cfg[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END cfg[23]
  PIN cfg[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 16.360 479.755 16.960 ;
    END
  END cfg[24]
  PIN cfg[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END cfg[25]
  PIN cfg[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END cfg[26]
  PIN cfg[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 325.770 486.475 326.050 490.475 ;
    END
  END cfg[27]
  PIN cfg[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 418.690 486.475 418.970 490.475 ;
    END
  END cfg[28]
  PIN cfg[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END cfg[29]
  PIN cfg[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END cfg[2]
  PIN cfg[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END cfg[30]
  PIN cfg[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 306.040 479.755 306.640 ;
    END
  END cfg[31]
  PIN cfg[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 452.730 486.475 453.010 490.475 ;
    END
  END cfg[32]
  PIN cfg[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.970 486.475 243.250 490.475 ;
    END
  END cfg[33]
  PIN cfg[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END cfg[34]
  PIN cfg[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END cfg[35]
  PIN cfg[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END cfg[36]
  PIN cfg[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END cfg[37]
  PIN cfg[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 53.080 479.755 53.680 ;
    END
  END cfg[38]
  PIN cfg[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 371.320 479.755 371.920 ;
    END
  END cfg[39]
  PIN cfg[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 443.400 479.755 444.000 ;
    END
  END cfg[3]
  PIN cfg[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END cfg[40]
  PIN cfg[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.050 486.475 81.330 490.475 ;
    END
  END cfg[41]
  PIN cfg[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END cfg[42]
  PIN cfg[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END cfg[43]
  PIN cfg[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 125.160 479.755 125.760 ;
    END
  END cfg[44]
  PIN cfg[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END cfg[45]
  PIN cfg[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 391.720 479.755 392.320 ;
    END
  END cfg[46]
  PIN cfg[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 384.650 486.475 384.930 490.475 ;
    END
  END cfg[47]
  PIN cfg[48]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END cfg[48]
  PIN cfg[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.450 486.475 76.730 490.475 ;
    END
  END cfg[49]
  PIN cfg[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 164.770 486.475 165.050 490.475 ;
    END
  END cfg[4]
  PIN cfg[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END cfg[50]
  PIN cfg[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.610 486.475 442.890 490.475 ;
    END
  END cfg[51]
  PIN cfg[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END cfg[52]
  PIN cfg[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END cfg[53]
  PIN cfg[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END cfg[54]
  PIN cfg[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END cfg[55]
  PIN cfg[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END cfg[56]
  PIN cfg[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END cfg[57]
  PIN cfg[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 369.930 486.475 370.210 490.475 ;
    END
  END cfg[58]
  PIN cfg[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END cfg[59]
  PIN cfg[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 374.530 486.475 374.810 490.475 ;
    END
  END cfg[5]
  PIN cfg[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 471.960 479.755 472.560 ;
    END
  END cfg[60]
  PIN cfg[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 284.280 479.755 284.880 ;
    END
  END cfg[61]
  PIN cfg[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 286.210 486.475 286.490 490.475 ;
    END
  END cfg[62]
  PIN cfg[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 140.120 479.755 140.720 ;
    END
  END cfg[63]
  PIN cfg[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END cfg[64]
  PIN cfg[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END cfg[65]
  PIN cfg[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.290 486.475 101.570 490.475 ;
    END
  END cfg[66]
  PIN cfg[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 486.475 3.130 490.475 ;
    END
  END cfg[67]
  PIN cfg[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END cfg[68]
  PIN cfg[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END cfg[69]
  PIN cfg[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 291.730 486.475 292.010 490.475 ;
    END
  END cfg[6]
  PIN cfg[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END cfg[70]
  PIN cfg[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 153.720 479.755 154.320 ;
    END
  END cfg[71]
  PIN cfg[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END cfg[72]
  PIN cfg[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END cfg[73]
  PIN cfg[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.250 486.475 159.530 490.475 ;
    END
  END cfg[74]
  PIN cfg[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END cfg[75]
  PIN cfg[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END cfg[76]
  PIN cfg[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END cfg[77]
  PIN cfg[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 31.320 479.755 31.920 ;
    END
  END cfg[78]
  PIN cfg[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.250 486.475 389.530 490.475 ;
    END
  END cfg[79]
  PIN cfg[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END cfg[7]
  PIN cfg[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END cfg[80]
  PIN cfg[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END cfg[81]
  PIN cfg[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END cfg[82]
  PIN cfg[83]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END cfg[83]
  PIN cfg[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 485.560 479.755 486.160 ;
    END
  END cfg[84]
  PIN cfg[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.090 486.475 345.370 490.475 ;
    END
  END cfg[85]
  PIN cfg[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 306.450 486.475 306.730 490.475 ;
    END
  END cfg[86]
  PIN cfg[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 190.440 479.755 191.040 ;
    END
  END cfg[87]
  PIN cfg[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 321.170 486.475 321.450 490.475 ;
    END
  END cfg[88]
  PIN cfg[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END cfg[89]
  PIN cfg[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 319.640 479.755 320.240 ;
    END
  END cfg[8]
  PIN cfg[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END cfg[90]
  PIN cfg[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END cfg[91]
  PIN cfg[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END cfg[92]
  PIN cfg[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END cfg[93]
  PIN cfg[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END cfg[94]
  PIN cfg[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 486.475 110.770 490.475 ;
    END
  END cfg[95]
  PIN cfg[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 96.600 479.755 97.200 ;
    END
  END cfg[96]
  PIN cfg[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END cfg[97]
  PIN cfg[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END cfg[98]
  PIN cfg[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END cfg[99]
  PIN cfg[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 399.880 479.755 400.480 ;
    END
  END cfg[9]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 457.330 486.475 457.610 490.475 ;
    END
  END clk
  PIN cset
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 475.755 219.000 479.755 219.600 ;
    END
  END cset
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 266.890 486.475 267.170 490.475 ;
    END
  END en
  PIN out0[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END out0[0]
  PIN out0[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 399.370 486.475 399.650 490.475 ;
    END
  END out0[10]
  PIN out0[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 255.720 479.755 256.320 ;
    END
  END out0[11]
  PIN out0[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 406.680 479.755 407.280 ;
    END
  END out0[12]
  PIN out0[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 291.080 479.755 291.680 ;
    END
  END out0[13]
  PIN out0[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 118.360 479.755 118.960 ;
    END
  END out0[14]
  PIN out0[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 173.970 486.475 174.250 490.475 ;
    END
  END out0[15]
  PIN out0[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 486.475 135.610 490.475 ;
    END
  END out0[16]
  PIN out0[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 486.475 120.890 490.475 ;
    END
  END out0[17]
  PIN out0[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END out0[18]
  PIN out0[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END out0[19]
  PIN out0[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 327.800 479.755 328.400 ;
    END
  END out0[1]
  PIN out0[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END out0[20]
  PIN out0[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END out0[21]
  PIN out0[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END out0[22]
  PIN out0[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END out0[23]
  PIN out0[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.530 486.475 213.810 490.475 ;
    END
  END out0[24]
  PIN out0[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.410 486.475 364.690 490.475 ;
    END
  END out0[25]
  PIN out0[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 384.920 479.755 385.520 ;
    END
  END out0[26]
  PIN out0[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 435.240 479.755 435.840 ;
    END
  END out0[27]
  PIN out0[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 486.475 51.890 490.475 ;
    END
  END out0[28]
  PIN out0[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 312.840 479.755 313.440 ;
    END
  END out0[29]
  PIN out0[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.010 486.475 438.290 490.475 ;
    END
  END out0[2]
  PIN out0[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END out0[30]
  PIN out0[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END out0[31]
  PIN out0[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END out0[3]
  PIN out0[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 38.120 479.755 38.720 ;
    END
  END out0[4]
  PIN out0[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 363.160 479.755 363.760 ;
    END
  END out0[5]
  PIN out0[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 330.370 486.475 330.650 490.475 ;
    END
  END out0[6]
  PIN out0[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 297.880 479.755 298.480 ;
    END
  END out0[7]
  PIN out0[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END out0[8]
  PIN out0[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 467.450 486.475 467.730 490.475 ;
    END
  END out0[9]
  PIN out1[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 315.650 486.475 315.930 490.475 ;
    END
  END out1[0]
  PIN out1[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 334.600 479.755 335.200 ;
    END
  END out1[10]
  PIN out1[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 421.640 479.755 422.240 ;
    END
  END out1[11]
  PIN out1[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END out1[12]
  PIN out1[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END out1[13]
  PIN out1[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.410 486.475 42.690 490.475 ;
    END
  END out1[14]
  PIN out1[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 296.330 486.475 296.610 490.475 ;
    END
  END out1[15]
  PIN out1[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END out1[16]
  PIN out1[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 182.280 479.755 182.880 ;
    END
  END out1[17]
  PIN out1[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 486.475 38.090 490.475 ;
    END
  END out1[18]
  PIN out1[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END out1[19]
  PIN out1[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END out1[1]
  PIN out1[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 457.000 479.755 457.600 ;
    END
  END out1[20]
  PIN out1[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 408.570 486.475 408.850 490.475 ;
    END
  END out1[21]
  PIN out1[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END out1[22]
  PIN out1[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END out1[23]
  PIN out1[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 125.210 486.475 125.490 490.475 ;
    END
  END out1[24]
  PIN out1[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END out1[25]
  PIN out1[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END out1[26]
  PIN out1[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 462.850 486.475 463.130 490.475 ;
    END
  END out1[27]
  PIN out1[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 161.880 479.755 162.480 ;
    END
  END out1[28]
  PIN out1[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END out1[29]
  PIN out1[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END out1[2]
  PIN out1[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END out1[30]
  PIN out1[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.970 486.475 13.250 490.475 ;
    END
  END out1[31]
  PIN out1[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 66.680 479.755 67.280 ;
    END
  END out1[3]
  PIN out1[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END out1[4]
  PIN out1[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END out1[5]
  PIN out1[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END out1[6]
  PIN out1[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 175.480 479.755 176.080 ;
    END
  END out1[7]
  PIN out1[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.010 486.475 208.290 490.475 ;
    END
  END out1[8]
  PIN out1[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 486.475 130.090 490.475 ;
    END
  END out1[9]
  PIN out2[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END out2[0]
  PIN out2[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END out2[10]
  PIN out2[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 486.475 96.050 490.475 ;
    END
  END out2[11]
  PIN out2[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 131.960 479.755 132.560 ;
    END
  END out2[12]
  PIN out2[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END out2[13]
  PIN out2[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END out2[14]
  PIN out2[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 237.450 486.475 237.730 490.475 ;
    END
  END out2[15]
  PIN out2[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 300.930 486.475 301.210 490.475 ;
    END
  END out2[16]
  PIN out2[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END out2[17]
  PIN out2[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 378.120 479.755 378.720 ;
    END
  END out2[18]
  PIN out2[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END out2[19]
  PIN out2[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END out2[1]
  PIN out2[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 144.530 486.475 144.810 490.475 ;
    END
  END out2[20]
  PIN out2[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END out2[21]
  PIN out2[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 478.760 479.755 479.360 ;
    END
  END out2[22]
  PIN out2[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END out2[23]
  PIN out2[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 225.800 479.755 226.400 ;
    END
  END out2[24]
  PIN out2[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END out2[25]
  PIN out2[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 46.280 479.755 46.880 ;
    END
  END out2[26]
  PIN out2[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END out2[27]
  PIN out2[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 427.890 486.475 428.170 490.475 ;
    END
  END out2[28]
  PIN out2[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END out2[29]
  PIN out2[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 232.850 486.475 233.130 490.475 ;
    END
  END out2[2]
  PIN out2[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END out2[30]
  PIN out2[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END out2[31]
  PIN out2[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.730 486.475 62.010 490.475 ;
    END
  END out2[3]
  PIN out2[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.130 486.475 379.410 490.475 ;
    END
  END out2[4]
  PIN out2[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 184.090 486.475 184.370 490.475 ;
    END
  END out2[5]
  PIN out2[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END out2[6]
  PIN out2[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 188.690 486.475 188.970 490.475 ;
    END
  END out2[7]
  PIN out2[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END out2[8]
  PIN out2[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 59.880 479.755 60.480 ;
    END
  END out2[9]
  PIN out3[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END out3[0]
  PIN out3[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.290 486.475 423.570 490.475 ;
    END
  END out3[10]
  PIN out3[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 271.490 486.475 271.770 490.475 ;
    END
  END out3[11]
  PIN out3[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 340.490 486.475 340.770 490.475 ;
    END
  END out3[12]
  PIN out3[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END out3[13]
  PIN out3[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END out3[14]
  PIN out3[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 276.120 479.755 276.720 ;
    END
  END out3[15]
  PIN out3[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END out3[16]
  PIN out3[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END out3[17]
  PIN out3[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 349.690 486.475 349.970 490.475 ;
    END
  END out3[18]
  PIN out3[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.170 486.475 91.450 490.475 ;
    END
  END out3[19]
  PIN out3[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 57.130 486.475 57.410 490.475 ;
    END
  END out3[1]
  PIN out3[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END out3[20]
  PIN out3[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END out3[21]
  PIN out3[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END out3[22]
  PIN out3[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 257.690 486.475 257.970 490.475 ;
    END
  END out3[23]
  PIN out3[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END out3[24]
  PIN out3[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 81.640 479.755 82.240 ;
    END
  END out3[25]
  PIN out3[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END out3[26]
  PIN out3[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 486.475 8.650 490.475 ;
    END
  END out3[27]
  PIN out3[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 355.210 486.475 355.490 490.475 ;
    END
  END out3[28]
  PIN out3[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 393.850 486.475 394.130 490.475 ;
    END
  END out3[29]
  PIN out3[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END out3[2]
  PIN out3[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END out3[30]
  PIN out3[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END out3[31]
  PIN out3[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END out3[3]
  PIN out3[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END out3[4]
  PIN out3[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.730 486.475 223.010 490.475 ;
    END
  END out3[5]
  PIN out3[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END out3[6]
  PIN out3[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 475.755 9.560 479.755 10.160 ;
    END
  END out3[7]
  PIN out3[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END out3[8]
  PIN out3[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 472.050 486.475 472.330 490.475 ;
    END
  END out3[9]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END rst
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 473.800 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 473.800 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.285 10.795 473.800 478.805 ;
      LAYER met1 ;
        RECT 2.830 6.840 476.950 486.160 ;
      LAYER met2 ;
        RECT 0.090 486.195 2.570 486.475 ;
        RECT 3.410 486.195 8.090 486.475 ;
        RECT 8.930 486.195 12.690 486.475 ;
        RECT 13.530 486.195 17.290 486.475 ;
        RECT 18.130 486.195 22.810 486.475 ;
        RECT 23.650 486.195 27.410 486.475 ;
        RECT 28.250 486.195 32.010 486.475 ;
        RECT 32.850 486.195 37.530 486.475 ;
        RECT 38.370 486.195 42.130 486.475 ;
        RECT 42.970 486.195 46.730 486.475 ;
        RECT 47.570 486.195 51.330 486.475 ;
        RECT 52.170 486.195 56.850 486.475 ;
        RECT 57.690 486.195 61.450 486.475 ;
        RECT 62.290 486.195 66.050 486.475 ;
        RECT 66.890 486.195 71.570 486.475 ;
        RECT 72.410 486.195 76.170 486.475 ;
        RECT 77.010 486.195 80.770 486.475 ;
        RECT 81.610 486.195 86.290 486.475 ;
        RECT 87.130 486.195 90.890 486.475 ;
        RECT 91.730 486.195 95.490 486.475 ;
        RECT 96.330 486.195 101.010 486.475 ;
        RECT 101.850 486.195 105.610 486.475 ;
        RECT 106.450 486.195 110.210 486.475 ;
        RECT 111.050 486.195 114.810 486.475 ;
        RECT 115.650 486.195 120.330 486.475 ;
        RECT 121.170 486.195 124.930 486.475 ;
        RECT 125.770 486.195 129.530 486.475 ;
        RECT 130.370 486.195 135.050 486.475 ;
        RECT 135.890 486.195 139.650 486.475 ;
        RECT 140.490 486.195 144.250 486.475 ;
        RECT 145.090 486.195 149.770 486.475 ;
        RECT 150.610 486.195 154.370 486.475 ;
        RECT 155.210 486.195 158.970 486.475 ;
        RECT 159.810 486.195 164.490 486.475 ;
        RECT 165.330 486.195 169.090 486.475 ;
        RECT 169.930 486.195 173.690 486.475 ;
        RECT 174.530 486.195 179.210 486.475 ;
        RECT 180.050 486.195 183.810 486.475 ;
        RECT 184.650 486.195 188.410 486.475 ;
        RECT 189.250 486.195 193.010 486.475 ;
        RECT 193.850 486.195 198.530 486.475 ;
        RECT 199.370 486.195 203.130 486.475 ;
        RECT 203.970 486.195 207.730 486.475 ;
        RECT 208.570 486.195 213.250 486.475 ;
        RECT 214.090 486.195 217.850 486.475 ;
        RECT 218.690 486.195 222.450 486.475 ;
        RECT 223.290 486.195 227.970 486.475 ;
        RECT 228.810 486.195 232.570 486.475 ;
        RECT 233.410 486.195 237.170 486.475 ;
        RECT 238.010 486.195 242.690 486.475 ;
        RECT 243.530 486.195 247.290 486.475 ;
        RECT 248.130 486.195 251.890 486.475 ;
        RECT 252.730 486.195 257.410 486.475 ;
        RECT 258.250 486.195 262.010 486.475 ;
        RECT 262.850 486.195 266.610 486.475 ;
        RECT 267.450 486.195 271.210 486.475 ;
        RECT 272.050 486.195 276.730 486.475 ;
        RECT 277.570 486.195 281.330 486.475 ;
        RECT 282.170 486.195 285.930 486.475 ;
        RECT 286.770 486.195 291.450 486.475 ;
        RECT 292.290 486.195 296.050 486.475 ;
        RECT 296.890 486.195 300.650 486.475 ;
        RECT 301.490 486.195 306.170 486.475 ;
        RECT 307.010 486.195 310.770 486.475 ;
        RECT 311.610 486.195 315.370 486.475 ;
        RECT 316.210 486.195 320.890 486.475 ;
        RECT 321.730 486.195 325.490 486.475 ;
        RECT 326.330 486.195 330.090 486.475 ;
        RECT 330.930 486.195 334.690 486.475 ;
        RECT 335.530 486.195 340.210 486.475 ;
        RECT 341.050 486.195 344.810 486.475 ;
        RECT 345.650 486.195 349.410 486.475 ;
        RECT 350.250 486.195 354.930 486.475 ;
        RECT 355.770 486.195 359.530 486.475 ;
        RECT 360.370 486.195 364.130 486.475 ;
        RECT 364.970 486.195 369.650 486.475 ;
        RECT 370.490 486.195 374.250 486.475 ;
        RECT 375.090 486.195 378.850 486.475 ;
        RECT 379.690 486.195 384.370 486.475 ;
        RECT 385.210 486.195 388.970 486.475 ;
        RECT 389.810 486.195 393.570 486.475 ;
        RECT 394.410 486.195 399.090 486.475 ;
        RECT 399.930 486.195 403.690 486.475 ;
        RECT 404.530 486.195 408.290 486.475 ;
        RECT 409.130 486.195 412.890 486.475 ;
        RECT 413.730 486.195 418.410 486.475 ;
        RECT 419.250 486.195 423.010 486.475 ;
        RECT 423.850 486.195 427.610 486.475 ;
        RECT 428.450 486.195 433.130 486.475 ;
        RECT 433.970 486.195 437.730 486.475 ;
        RECT 438.570 486.195 442.330 486.475 ;
        RECT 443.170 486.195 447.850 486.475 ;
        RECT 448.690 486.195 452.450 486.475 ;
        RECT 453.290 486.195 457.050 486.475 ;
        RECT 457.890 486.195 462.570 486.475 ;
        RECT 463.410 486.195 467.170 486.475 ;
        RECT 468.010 486.195 471.770 486.475 ;
        RECT 472.610 486.195 476.920 486.475 ;
        RECT 0.090 4.280 476.920 486.195 ;
        RECT 0.090 4.000 2.570 4.280 ;
        RECT 3.410 4.000 7.170 4.280 ;
        RECT 8.010 4.000 11.770 4.280 ;
        RECT 12.610 4.000 16.370 4.280 ;
        RECT 17.210 4.000 21.890 4.280 ;
        RECT 22.730 4.000 26.490 4.280 ;
        RECT 27.330 4.000 31.090 4.280 ;
        RECT 31.930 4.000 36.610 4.280 ;
        RECT 37.450 4.000 41.210 4.280 ;
        RECT 42.050 4.000 45.810 4.280 ;
        RECT 46.650 4.000 51.330 4.280 ;
        RECT 52.170 4.000 55.930 4.280 ;
        RECT 56.770 4.000 60.530 4.280 ;
        RECT 61.370 4.000 66.050 4.280 ;
        RECT 66.890 4.000 70.650 4.280 ;
        RECT 71.490 4.000 75.250 4.280 ;
        RECT 76.090 4.000 79.850 4.280 ;
        RECT 80.690 4.000 85.370 4.280 ;
        RECT 86.210 4.000 89.970 4.280 ;
        RECT 90.810 4.000 94.570 4.280 ;
        RECT 95.410 4.000 100.090 4.280 ;
        RECT 100.930 4.000 104.690 4.280 ;
        RECT 105.530 4.000 109.290 4.280 ;
        RECT 110.130 4.000 114.810 4.280 ;
        RECT 115.650 4.000 119.410 4.280 ;
        RECT 120.250 4.000 124.010 4.280 ;
        RECT 124.850 4.000 129.530 4.280 ;
        RECT 130.370 4.000 134.130 4.280 ;
        RECT 134.970 4.000 138.730 4.280 ;
        RECT 139.570 4.000 144.250 4.280 ;
        RECT 145.090 4.000 148.850 4.280 ;
        RECT 149.690 4.000 153.450 4.280 ;
        RECT 154.290 4.000 158.050 4.280 ;
        RECT 158.890 4.000 163.570 4.280 ;
        RECT 164.410 4.000 168.170 4.280 ;
        RECT 169.010 4.000 172.770 4.280 ;
        RECT 173.610 4.000 178.290 4.280 ;
        RECT 179.130 4.000 182.890 4.280 ;
        RECT 183.730 4.000 187.490 4.280 ;
        RECT 188.330 4.000 193.010 4.280 ;
        RECT 193.850 4.000 197.610 4.280 ;
        RECT 198.450 4.000 202.210 4.280 ;
        RECT 203.050 4.000 207.730 4.280 ;
        RECT 208.570 4.000 212.330 4.280 ;
        RECT 213.170 4.000 216.930 4.280 ;
        RECT 217.770 4.000 221.530 4.280 ;
        RECT 222.370 4.000 227.050 4.280 ;
        RECT 227.890 4.000 231.650 4.280 ;
        RECT 232.490 4.000 236.250 4.280 ;
        RECT 237.090 4.000 241.770 4.280 ;
        RECT 242.610 4.000 246.370 4.280 ;
        RECT 247.210 4.000 250.970 4.280 ;
        RECT 251.810 4.000 256.490 4.280 ;
        RECT 257.330 4.000 261.090 4.280 ;
        RECT 261.930 4.000 265.690 4.280 ;
        RECT 266.530 4.000 271.210 4.280 ;
        RECT 272.050 4.000 275.810 4.280 ;
        RECT 276.650 4.000 280.410 4.280 ;
        RECT 281.250 4.000 285.930 4.280 ;
        RECT 286.770 4.000 290.530 4.280 ;
        RECT 291.370 4.000 295.130 4.280 ;
        RECT 295.970 4.000 299.730 4.280 ;
        RECT 300.570 4.000 305.250 4.280 ;
        RECT 306.090 4.000 309.850 4.280 ;
        RECT 310.690 4.000 314.450 4.280 ;
        RECT 315.290 4.000 319.970 4.280 ;
        RECT 320.810 4.000 324.570 4.280 ;
        RECT 325.410 4.000 329.170 4.280 ;
        RECT 330.010 4.000 334.690 4.280 ;
        RECT 335.530 4.000 339.290 4.280 ;
        RECT 340.130 4.000 343.890 4.280 ;
        RECT 344.730 4.000 349.410 4.280 ;
        RECT 350.250 4.000 354.010 4.280 ;
        RECT 354.850 4.000 358.610 4.280 ;
        RECT 359.450 4.000 364.130 4.280 ;
        RECT 364.970 4.000 368.730 4.280 ;
        RECT 369.570 4.000 373.330 4.280 ;
        RECT 374.170 4.000 377.930 4.280 ;
        RECT 378.770 4.000 383.450 4.280 ;
        RECT 384.290 4.000 388.050 4.280 ;
        RECT 388.890 4.000 392.650 4.280 ;
        RECT 393.490 4.000 398.170 4.280 ;
        RECT 399.010 4.000 402.770 4.280 ;
        RECT 403.610 4.000 407.370 4.280 ;
        RECT 408.210 4.000 412.890 4.280 ;
        RECT 413.730 4.000 417.490 4.280 ;
        RECT 418.330 4.000 422.090 4.280 ;
        RECT 422.930 4.000 427.610 4.280 ;
        RECT 428.450 4.000 432.210 4.280 ;
        RECT 433.050 4.000 436.810 4.280 ;
        RECT 437.650 4.000 441.410 4.280 ;
        RECT 442.250 4.000 446.930 4.280 ;
        RECT 447.770 4.000 451.530 4.280 ;
        RECT 452.370 4.000 456.130 4.280 ;
        RECT 456.970 4.000 461.650 4.280 ;
        RECT 462.490 4.000 466.250 4.280 ;
        RECT 467.090 4.000 470.850 4.280 ;
        RECT 471.690 4.000 476.370 4.280 ;
      LAYER met3 ;
        RECT 0.065 485.160 475.355 486.025 ;
        RECT 0.065 481.120 475.755 485.160 ;
        RECT 4.400 479.760 475.755 481.120 ;
        RECT 4.400 479.720 475.355 479.760 ;
        RECT 0.065 478.360 475.355 479.720 ;
        RECT 0.065 474.320 475.755 478.360 ;
        RECT 4.400 472.960 475.755 474.320 ;
        RECT 4.400 472.920 475.355 472.960 ;
        RECT 0.065 471.560 475.355 472.920 ;
        RECT 0.065 466.160 475.755 471.560 ;
        RECT 4.400 464.760 475.355 466.160 ;
        RECT 0.065 459.360 475.755 464.760 ;
        RECT 4.400 458.000 475.755 459.360 ;
        RECT 4.400 457.960 475.355 458.000 ;
        RECT 0.065 456.600 475.355 457.960 ;
        RECT 0.065 452.560 475.755 456.600 ;
        RECT 4.400 451.200 475.755 452.560 ;
        RECT 4.400 451.160 475.355 451.200 ;
        RECT 0.065 449.800 475.355 451.160 ;
        RECT 0.065 444.400 475.755 449.800 ;
        RECT 4.400 443.000 475.355 444.400 ;
        RECT 0.065 437.600 475.755 443.000 ;
        RECT 4.400 436.240 475.755 437.600 ;
        RECT 4.400 436.200 475.355 436.240 ;
        RECT 0.065 434.840 475.355 436.200 ;
        RECT 0.065 430.800 475.755 434.840 ;
        RECT 4.400 429.440 475.755 430.800 ;
        RECT 4.400 429.400 475.355 429.440 ;
        RECT 0.065 428.040 475.355 429.400 ;
        RECT 0.065 424.000 475.755 428.040 ;
        RECT 4.400 422.640 475.755 424.000 ;
        RECT 4.400 422.600 475.355 422.640 ;
        RECT 0.065 421.240 475.355 422.600 ;
        RECT 0.065 415.840 475.755 421.240 ;
        RECT 4.400 414.480 475.755 415.840 ;
        RECT 4.400 414.440 475.355 414.480 ;
        RECT 0.065 413.080 475.355 414.440 ;
        RECT 0.065 409.040 475.755 413.080 ;
        RECT 4.400 407.680 475.755 409.040 ;
        RECT 4.400 407.640 475.355 407.680 ;
        RECT 0.065 406.280 475.355 407.640 ;
        RECT 0.065 402.240 475.755 406.280 ;
        RECT 4.400 400.880 475.755 402.240 ;
        RECT 4.400 400.840 475.355 400.880 ;
        RECT 0.065 399.480 475.355 400.840 ;
        RECT 0.065 394.080 475.755 399.480 ;
        RECT 4.400 392.720 475.755 394.080 ;
        RECT 4.400 392.680 475.355 392.720 ;
        RECT 0.065 391.320 475.355 392.680 ;
        RECT 0.065 387.280 475.755 391.320 ;
        RECT 4.400 385.920 475.755 387.280 ;
        RECT 4.400 385.880 475.355 385.920 ;
        RECT 0.065 384.520 475.355 385.880 ;
        RECT 0.065 380.480 475.755 384.520 ;
        RECT 4.400 379.120 475.755 380.480 ;
        RECT 4.400 379.080 475.355 379.120 ;
        RECT 0.065 377.720 475.355 379.080 ;
        RECT 0.065 372.320 475.755 377.720 ;
        RECT 4.400 370.920 475.355 372.320 ;
        RECT 0.065 365.520 475.755 370.920 ;
        RECT 4.400 364.160 475.755 365.520 ;
        RECT 4.400 364.120 475.355 364.160 ;
        RECT 0.065 362.760 475.355 364.120 ;
        RECT 0.065 358.720 475.755 362.760 ;
        RECT 4.400 357.360 475.755 358.720 ;
        RECT 4.400 357.320 475.355 357.360 ;
        RECT 0.065 355.960 475.355 357.320 ;
        RECT 0.065 350.560 475.755 355.960 ;
        RECT 4.400 349.160 475.355 350.560 ;
        RECT 0.065 343.760 475.755 349.160 ;
        RECT 4.400 342.400 475.755 343.760 ;
        RECT 4.400 342.360 475.355 342.400 ;
        RECT 0.065 341.000 475.355 342.360 ;
        RECT 0.065 336.960 475.755 341.000 ;
        RECT 4.400 335.600 475.755 336.960 ;
        RECT 4.400 335.560 475.355 335.600 ;
        RECT 0.065 334.200 475.355 335.560 ;
        RECT 0.065 328.800 475.755 334.200 ;
        RECT 4.400 327.400 475.355 328.800 ;
        RECT 0.065 322.000 475.755 327.400 ;
        RECT 4.400 320.640 475.755 322.000 ;
        RECT 4.400 320.600 475.355 320.640 ;
        RECT 0.065 319.240 475.355 320.600 ;
        RECT 0.065 315.200 475.755 319.240 ;
        RECT 4.400 313.840 475.755 315.200 ;
        RECT 4.400 313.800 475.355 313.840 ;
        RECT 0.065 312.440 475.355 313.800 ;
        RECT 0.065 308.400 475.755 312.440 ;
        RECT 4.400 307.040 475.755 308.400 ;
        RECT 4.400 307.000 475.355 307.040 ;
        RECT 0.065 305.640 475.355 307.000 ;
        RECT 0.065 300.240 475.755 305.640 ;
        RECT 4.400 298.880 475.755 300.240 ;
        RECT 4.400 298.840 475.355 298.880 ;
        RECT 0.065 297.480 475.355 298.840 ;
        RECT 0.065 293.440 475.755 297.480 ;
        RECT 4.400 292.080 475.755 293.440 ;
        RECT 4.400 292.040 475.355 292.080 ;
        RECT 0.065 290.680 475.355 292.040 ;
        RECT 0.065 286.640 475.755 290.680 ;
        RECT 4.400 285.280 475.755 286.640 ;
        RECT 4.400 285.240 475.355 285.280 ;
        RECT 0.065 283.880 475.355 285.240 ;
        RECT 0.065 278.480 475.755 283.880 ;
        RECT 4.400 277.120 475.755 278.480 ;
        RECT 4.400 277.080 475.355 277.120 ;
        RECT 0.065 275.720 475.355 277.080 ;
        RECT 0.065 271.680 475.755 275.720 ;
        RECT 4.400 270.320 475.755 271.680 ;
        RECT 4.400 270.280 475.355 270.320 ;
        RECT 0.065 268.920 475.355 270.280 ;
        RECT 0.065 264.880 475.755 268.920 ;
        RECT 4.400 263.520 475.755 264.880 ;
        RECT 4.400 263.480 475.355 263.520 ;
        RECT 0.065 262.120 475.355 263.480 ;
        RECT 0.065 256.720 475.755 262.120 ;
        RECT 4.400 255.320 475.355 256.720 ;
        RECT 0.065 249.920 475.755 255.320 ;
        RECT 4.400 248.560 475.755 249.920 ;
        RECT 4.400 248.520 475.355 248.560 ;
        RECT 0.065 247.160 475.355 248.520 ;
        RECT 0.065 243.120 475.755 247.160 ;
        RECT 4.400 241.760 475.755 243.120 ;
        RECT 4.400 241.720 475.355 241.760 ;
        RECT 0.065 240.360 475.355 241.720 ;
        RECT 0.065 234.960 475.755 240.360 ;
        RECT 4.400 233.560 475.355 234.960 ;
        RECT 0.065 228.160 475.755 233.560 ;
        RECT 4.400 226.800 475.755 228.160 ;
        RECT 4.400 226.760 475.355 226.800 ;
        RECT 0.065 225.400 475.355 226.760 ;
        RECT 0.065 221.360 475.755 225.400 ;
        RECT 4.400 220.000 475.755 221.360 ;
        RECT 4.400 219.960 475.355 220.000 ;
        RECT 0.065 218.600 475.355 219.960 ;
        RECT 0.065 214.560 475.755 218.600 ;
        RECT 4.400 213.200 475.755 214.560 ;
        RECT 4.400 213.160 475.355 213.200 ;
        RECT 0.065 211.800 475.355 213.160 ;
        RECT 0.065 206.400 475.755 211.800 ;
        RECT 4.400 205.040 475.755 206.400 ;
        RECT 4.400 205.000 475.355 205.040 ;
        RECT 0.065 203.640 475.355 205.000 ;
        RECT 0.065 199.600 475.755 203.640 ;
        RECT 4.400 198.240 475.755 199.600 ;
        RECT 4.400 198.200 475.355 198.240 ;
        RECT 0.065 196.840 475.355 198.200 ;
        RECT 0.065 192.800 475.755 196.840 ;
        RECT 4.400 191.440 475.755 192.800 ;
        RECT 4.400 191.400 475.355 191.440 ;
        RECT 0.065 190.040 475.355 191.400 ;
        RECT 0.065 184.640 475.755 190.040 ;
        RECT 4.400 183.280 475.755 184.640 ;
        RECT 4.400 183.240 475.355 183.280 ;
        RECT 0.065 181.880 475.355 183.240 ;
        RECT 0.065 177.840 475.755 181.880 ;
        RECT 4.400 176.480 475.755 177.840 ;
        RECT 4.400 176.440 475.355 176.480 ;
        RECT 0.065 175.080 475.355 176.440 ;
        RECT 0.065 171.040 475.755 175.080 ;
        RECT 4.400 169.680 475.755 171.040 ;
        RECT 4.400 169.640 475.355 169.680 ;
        RECT 0.065 168.280 475.355 169.640 ;
        RECT 0.065 162.880 475.755 168.280 ;
        RECT 4.400 161.480 475.355 162.880 ;
        RECT 0.065 156.080 475.755 161.480 ;
        RECT 4.400 154.720 475.755 156.080 ;
        RECT 4.400 154.680 475.355 154.720 ;
        RECT 0.065 153.320 475.355 154.680 ;
        RECT 0.065 149.280 475.755 153.320 ;
        RECT 4.400 147.920 475.755 149.280 ;
        RECT 4.400 147.880 475.355 147.920 ;
        RECT 0.065 146.520 475.355 147.880 ;
        RECT 0.065 141.120 475.755 146.520 ;
        RECT 4.400 139.720 475.355 141.120 ;
        RECT 0.065 134.320 475.755 139.720 ;
        RECT 4.400 132.960 475.755 134.320 ;
        RECT 4.400 132.920 475.355 132.960 ;
        RECT 0.065 131.560 475.355 132.920 ;
        RECT 0.065 127.520 475.755 131.560 ;
        RECT 4.400 126.160 475.755 127.520 ;
        RECT 4.400 126.120 475.355 126.160 ;
        RECT 0.065 124.760 475.355 126.120 ;
        RECT 0.065 119.360 475.755 124.760 ;
        RECT 4.400 117.960 475.355 119.360 ;
        RECT 0.065 112.560 475.755 117.960 ;
        RECT 4.400 111.200 475.755 112.560 ;
        RECT 4.400 111.160 475.355 111.200 ;
        RECT 0.065 109.800 475.355 111.160 ;
        RECT 0.065 105.760 475.755 109.800 ;
        RECT 4.400 104.400 475.755 105.760 ;
        RECT 4.400 104.360 475.355 104.400 ;
        RECT 0.065 103.000 475.355 104.360 ;
        RECT 0.065 98.960 475.755 103.000 ;
        RECT 4.400 97.600 475.755 98.960 ;
        RECT 4.400 97.560 475.355 97.600 ;
        RECT 0.065 96.200 475.355 97.560 ;
        RECT 0.065 90.800 475.755 96.200 ;
        RECT 4.400 89.440 475.755 90.800 ;
        RECT 4.400 89.400 475.355 89.440 ;
        RECT 0.065 88.040 475.355 89.400 ;
        RECT 0.065 84.000 475.755 88.040 ;
        RECT 4.400 82.640 475.755 84.000 ;
        RECT 4.400 82.600 475.355 82.640 ;
        RECT 0.065 81.240 475.355 82.600 ;
        RECT 0.065 77.200 475.755 81.240 ;
        RECT 4.400 75.840 475.755 77.200 ;
        RECT 4.400 75.800 475.355 75.840 ;
        RECT 0.065 74.440 475.355 75.800 ;
        RECT 0.065 69.040 475.755 74.440 ;
        RECT 4.400 67.680 475.755 69.040 ;
        RECT 4.400 67.640 475.355 67.680 ;
        RECT 0.065 66.280 475.355 67.640 ;
        RECT 0.065 62.240 475.755 66.280 ;
        RECT 4.400 60.880 475.755 62.240 ;
        RECT 4.400 60.840 475.355 60.880 ;
        RECT 0.065 59.480 475.355 60.840 ;
        RECT 0.065 55.440 475.755 59.480 ;
        RECT 4.400 54.080 475.755 55.440 ;
        RECT 4.400 54.040 475.355 54.080 ;
        RECT 0.065 52.680 475.355 54.040 ;
        RECT 0.065 47.280 475.755 52.680 ;
        RECT 4.400 45.880 475.355 47.280 ;
        RECT 0.065 40.480 475.755 45.880 ;
        RECT 4.400 39.120 475.755 40.480 ;
        RECT 4.400 39.080 475.355 39.120 ;
        RECT 0.065 37.720 475.355 39.080 ;
        RECT 0.065 33.680 475.755 37.720 ;
        RECT 4.400 32.320 475.755 33.680 ;
        RECT 4.400 32.280 475.355 32.320 ;
        RECT 0.065 30.920 475.355 32.280 ;
        RECT 0.065 25.520 475.755 30.920 ;
        RECT 4.400 24.120 475.355 25.520 ;
        RECT 0.065 18.720 475.755 24.120 ;
        RECT 4.400 17.360 475.755 18.720 ;
        RECT 4.400 17.320 475.355 17.360 ;
        RECT 0.065 15.960 475.355 17.320 ;
        RECT 0.065 11.920 475.755 15.960 ;
        RECT 4.400 10.560 475.755 11.920 ;
        RECT 4.400 10.520 475.355 10.560 ;
        RECT 0.065 9.160 475.355 10.520 ;
        RECT 0.065 4.255 475.755 9.160 ;
      LAYER met4 ;
        RECT 9.495 10.640 434.865 478.960 ;
      LAYER met5 ;
        RECT 5.520 179.670 473.800 411.040 ;
  END
END mac_cluster
END LIBRARY

