VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mac_cluster
  CLASS BLOCK ;
  FOREIGN mac_cluster ;
  ORIGIN 0.000 0.000 ;
  SIZE 510.265 BY 520.985 ;
  PIN A0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.530 516.985 190.810 520.985 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 277.480 510.265 278.080 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 429.730 516.985 430.010 520.985 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.170 516.985 206.450 520.985 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END A0[7]
  PIN A1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.410 516.985 180.690 520.985 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 477.400 510.265 478.000 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 268.730 516.985 269.010 520.985 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 294.490 516.985 294.770 520.985 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 516.985 19.690 520.985 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 278.850 516.985 279.130 520.985 ;
    END
  END A1[7]
  PIN A2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.010 516.985 461.290 520.985 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END A2[6]
  PIN A2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 454.280 510.265 454.880 ;
    END
  END A2[7]
  PIN A3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.970 516.985 243.250 520.985 ;
    END
  END A3[0]
  PIN A3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END A3[1]
  PIN A3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 476.650 516.985 476.930 520.985 ;
    END
  END A3[2]
  PIN A3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 211.690 516.985 211.970 520.985 ;
    END
  END A3[3]
  PIN A3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END A3[4]
  PIN A3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END A3[5]
  PIN A3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END A3[6]
  PIN A3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.930 516.985 71.210 520.985 ;
    END
  END A3[7]
  PIN B0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END B0[0]
  PIN B0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END B0[1]
  PIN B0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END B0[2]
  PIN B0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END B0[3]
  PIN B0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 224.440 510.265 225.040 ;
    END
  END B0[4]
  PIN B0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.930 516.985 232.210 520.985 ;
    END
  END B0[5]
  PIN B0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.450 516.985 76.730 520.985 ;
    END
  END B0[6]
  PIN B0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END B0[7]
  PIN B1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.130 516.985 149.410 520.985 ;
    END
  END B1[0]
  PIN B1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 378.120 510.265 378.720 ;
    END
  END B1[1]
  PIN B1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 155.080 510.265 155.680 ;
    END
  END B1[2]
  PIN B1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END B1[3]
  PIN B1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 382.810 516.985 383.090 520.985 ;
    END
  END B1[4]
  PIN B1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END B1[5]
  PIN B1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.250 516.985 159.530 520.985 ;
    END
  END B1[6]
  PIN B1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 247.560 510.265 248.160 ;
    END
  END B1[7]
  PIN B2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END B2[0]
  PIN B2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END B2[1]
  PIN B2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END B2[2]
  PIN B2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 117.000 510.265 117.600 ;
    END
  END B2[3]
  PIN B2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 164.770 516.985 165.050 520.985 ;
    END
  END B2[4]
  PIN B2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 516.985 24.290 520.985 ;
    END
  END B2[5]
  PIN B2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END B2[6]
  PIN B2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 285.640 510.265 286.240 ;
    END
  END B2[7]
  PIN B3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 78.920 510.265 79.520 ;
    END
  END B3[0]
  PIN B3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END B3[1]
  PIN B3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END B3[2]
  PIN B3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 493.720 510.265 494.320 ;
    END
  END B3[3]
  PIN B3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 216.280 510.265 216.880 ;
    END
  END B3[4]
  PIN B3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 516.985 29.810 520.985 ;
    END
  END B3[5]
  PIN B3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END B3[6]
  PIN B3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 108.840 510.265 109.440 ;
    END
  END B3[7]
  PIN cfg[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.210 516.985 263.490 520.985 ;
    END
  END cfg[0]
  PIN cfg[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END cfg[100]
  PIN cfg[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END cfg[101]
  PIN cfg[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END cfg[102]
  PIN cfg[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 516.985 50.970 520.985 ;
    END
  END cfg[103]
  PIN cfg[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END cfg[104]
  PIN cfg[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END cfg[105]
  PIN cfg[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 439.320 510.265 439.920 ;
    END
  END cfg[106]
  PIN cfg[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END cfg[107]
  PIN cfg[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END cfg[108]
  PIN cfg[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.330 516.985 112.610 520.985 ;
    END
  END cfg[109]
  PIN cfg[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END cfg[10]
  PIN cfg[110]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END cfg[110]
  PIN cfg[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END cfg[111]
  PIN cfg[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END cfg[112]
  PIN cfg[113]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 209.480 510.265 210.080 ;
    END
  END cfg[113]
  PIN cfg[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 255.720 510.265 256.320 ;
    END
  END cfg[114]
  PIN cfg[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.090 516.985 92.370 520.985 ;
    END
  END cfg[115]
  PIN cfg[116]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END cfg[116]
  PIN cfg[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 439.850 516.985 440.130 520.985 ;
    END
  END cfg[117]
  PIN cfg[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END cfg[118]
  PIN cfg[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END cfg[119]
  PIN cfg[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END cfg[11]
  PIN cfg[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.370 516.985 123.650 520.985 ;
    END
  END cfg[120]
  PIN cfg[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 24.520 510.265 25.120 ;
    END
  END cfg[121]
  PIN cfg[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END cfg[122]
  PIN cfg[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END cfg[123]
  PIN cfg[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 369.960 510.265 370.560 ;
    END
  END cfg[124]
  PIN cfg[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 516.985 35.330 520.985 ;
    END
  END cfg[125]
  PIN cfg[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 262.520 510.265 263.120 ;
    END
  END cfg[126]
  PIN cfg[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END cfg[127]
  PIN cfg[128]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END cfg[128]
  PIN cfg[129]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END cfg[129]
  PIN cfg[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END cfg[12]
  PIN cfg[130]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END cfg[130]
  PIN cfg[131]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.050 516.985 357.330 520.985 ;
    END
  END cfg[131]
  PIN cfg[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 331.290 516.985 331.570 520.985 ;
    END
  END cfg[13]
  PIN cfg[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END cfg[14]
  PIN cfg[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END cfg[15]
  PIN cfg[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END cfg[16]
  PIN cfg[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.010 516.985 300.290 520.985 ;
    END
  END cfg[17]
  PIN cfg[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 363.160 510.265 363.760 ;
    END
  END cfg[18]
  PIN cfg[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END cfg[19]
  PIN cfg[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END cfg[1]
  PIN cfg[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 216.290 516.985 216.570 520.985 ;
    END
  END cfg[20]
  PIN cfg[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 93.880 510.265 94.480 ;
    END
  END cfg[21]
  PIN cfg[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 178.200 510.265 178.800 ;
    END
  END cfg[22]
  PIN cfg[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END cfg[23]
  PIN cfg[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 16.360 510.265 16.960 ;
    END
  END cfg[24]
  PIN cfg[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 501.490 0.000 501.770 4.000 ;
    END
  END cfg[25]
  PIN cfg[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END cfg[26]
  PIN cfg[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 346.010 516.985 346.290 520.985 ;
    END
  END cfg[27]
  PIN cfg[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 445.370 516.985 445.650 520.985 ;
    END
  END cfg[28]
  PIN cfg[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END cfg[29]
  PIN cfg[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END cfg[2]
  PIN cfg[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END cfg[30]
  PIN cfg[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 323.720 510.265 324.320 ;
    END
  END cfg[31]
  PIN cfg[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 481.250 516.985 481.530 520.985 ;
    END
  END cfg[32]
  PIN cfg[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 257.690 516.985 257.970 520.985 ;
    END
  END cfg[33]
  PIN cfg[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END cfg[34]
  PIN cfg[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END cfg[35]
  PIN cfg[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END cfg[36]
  PIN cfg[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END cfg[37]
  PIN cfg[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 55.800 510.265 56.400 ;
    END
  END cfg[38]
  PIN cfg[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 393.080 510.265 393.680 ;
    END
  END cfg[39]
  PIN cfg[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 470.600 510.265 471.200 ;
    END
  END cfg[3]
  PIN cfg[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END cfg[40]
  PIN cfg[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.570 516.985 86.850 520.985 ;
    END
  END cfg[41]
  PIN cfg[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END cfg[42]
  PIN cfg[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END cfg[43]
  PIN cfg[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 131.960 510.265 132.560 ;
    END
  END cfg[44]
  PIN cfg[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END cfg[45]
  PIN cfg[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 416.200 510.265 416.800 ;
    END
  END cfg[46]
  PIN cfg[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.570 516.985 408.850 520.985 ;
    END
  END cfg[47]
  PIN cfg[48]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END cfg[48]
  PIN cfg[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.050 516.985 81.330 520.985 ;
    END
  END cfg[49]
  PIN cfg[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.890 516.985 175.170 520.985 ;
    END
  END cfg[4]
  PIN cfg[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END cfg[50]
  PIN cfg[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.130 516.985 471.410 520.985 ;
    END
  END cfg[51]
  PIN cfg[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END cfg[52]
  PIN cfg[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END cfg[53]
  PIN cfg[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END cfg[54]
  PIN cfg[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END cfg[55]
  PIN cfg[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END cfg[56]
  PIN cfg[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END cfg[57]
  PIN cfg[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.930 516.985 393.210 520.985 ;
    END
  END cfg[58]
  PIN cfg[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END cfg[59]
  PIN cfg[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 398.450 516.985 398.730 520.985 ;
    END
  END cfg[5]
  PIN cfg[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 500.520 510.265 501.120 ;
    END
  END cfg[60]
  PIN cfg[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 300.600 510.265 301.200 ;
    END
  END cfg[61]
  PIN cfg[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 304.610 516.985 304.890 520.985 ;
    END
  END cfg[62]
  PIN cfg[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 146.920 510.265 147.520 ;
    END
  END cfg[63]
  PIN cfg[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END cfg[64]
  PIN cfg[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END cfg[65]
  PIN cfg[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 107.730 516.985 108.010 520.985 ;
    END
  END cfg[66]
  PIN cfg[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 516.985 4.050 520.985 ;
    END
  END cfg[67]
  PIN cfg[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 480.330 0.000 480.610 4.000 ;
    END
  END cfg[68]
  PIN cfg[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END cfg[69]
  PIN cfg[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 310.130 516.985 310.410 520.985 ;
    END
  END cfg[6]
  PIN cfg[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END cfg[70]
  PIN cfg[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 163.240 510.265 163.840 ;
    END
  END cfg[71]
  PIN cfg[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END cfg[72]
  PIN cfg[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END cfg[73]
  PIN cfg[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.370 516.985 169.650 520.985 ;
    END
  END cfg[74]
  PIN cfg[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END cfg[75]
  PIN cfg[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END cfg[76]
  PIN cfg[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END cfg[77]
  PIN cfg[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 32.680 510.265 33.280 ;
    END
  END cfg[78]
  PIN cfg[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.090 516.985 414.370 520.985 ;
    END
  END cfg[79]
  PIN cfg[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END cfg[7]
  PIN cfg[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END cfg[80]
  PIN cfg[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END cfg[81]
  PIN cfg[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END cfg[82]
  PIN cfg[83]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END cfg[83]
  PIN cfg[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.010 516.985 507.290 520.985 ;
    END
  END cfg[84]
  PIN cfg[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 367.170 516.985 367.450 520.985 ;
    END
  END cfg[85]
  PIN cfg[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 325.770 516.985 326.050 520.985 ;
    END
  END cfg[86]
  PIN cfg[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 201.320 510.265 201.920 ;
    END
  END cfg[87]
  PIN cfg[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 341.410 516.985 341.690 520.985 ;
    END
  END cfg[88]
  PIN cfg[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END cfg[89]
  PIN cfg[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 340.040 510.265 340.640 ;
    END
  END cfg[8]
  PIN cfg[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END cfg[90]
  PIN cfg[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END cfg[91]
  PIN cfg[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END cfg[92]
  PIN cfg[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END cfg[93]
  PIN cfg[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END cfg[94]
  PIN cfg[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.850 516.985 118.130 520.985 ;
    END
  END cfg[95]
  PIN cfg[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 102.040 510.265 102.640 ;
    END
  END cfg[96]
  PIN cfg[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END cfg[97]
  PIN cfg[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END cfg[98]
  PIN cfg[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END cfg[99]
  PIN cfg[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 424.360 510.265 424.960 ;
    END
  END cfg[9]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 486.770 516.985 487.050 520.985 ;
    END
  END clk
  PIN cset
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 506.265 232.600 510.265 233.200 ;
    END
  END cset
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 284.370 516.985 284.650 520.985 ;
    END
  END en
  PIN out0[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END out0[0]
  PIN out0[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 424.210 516.985 424.490 520.985 ;
    END
  END out0[10]
  PIN out0[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 270.680 510.265 271.280 ;
    END
  END out0[11]
  PIN out0[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 431.160 510.265 431.760 ;
    END
  END out0[12]
  PIN out0[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 308.760 510.265 309.360 ;
    END
  END out0[13]
  PIN out0[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 125.160 510.265 125.760 ;
    END
  END out0[14]
  PIN out0[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.010 516.985 185.290 520.985 ;
    END
  END out0[15]
  PIN out0[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 143.610 516.985 143.890 520.985 ;
    END
  END out0[16]
  PIN out0[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.970 516.985 128.250 520.985 ;
    END
  END out0[17]
  PIN out0[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END out0[18]
  PIN out0[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END out0[19]
  PIN out0[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 346.840 510.265 347.440 ;
    END
  END out0[1]
  PIN out0[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END out0[20]
  PIN out0[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END out0[21]
  PIN out0[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END out0[22]
  PIN out0[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END out0[23]
  PIN out0[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 227.330 516.985 227.610 520.985 ;
    END
  END out0[24]
  PIN out0[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.330 516.985 388.610 520.985 ;
    END
  END out0[25]
  PIN out0[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 408.040 510.265 408.640 ;
    END
  END out0[26]
  PIN out0[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 462.440 510.265 463.040 ;
    END
  END out0[27]
  PIN out0[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 516.985 55.570 520.985 ;
    END
  END out0[28]
  PIN out0[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 331.880 510.265 332.480 ;
    END
  END out0[29]
  PIN out0[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 465.610 516.985 465.890 520.985 ;
    END
  END out0[2]
  PIN out0[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END out0[30]
  PIN out0[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END out0[31]
  PIN out0[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END out0[3]
  PIN out0[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 39.480 510.265 40.080 ;
    END
  END out0[4]
  PIN out0[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 386.280 510.265 386.880 ;
    END
  END out0[5]
  PIN out0[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 351.530 516.985 351.810 520.985 ;
    END
  END out0[6]
  PIN out0[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 316.920 510.265 317.520 ;
    END
  END out0[7]
  PIN out0[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END out0[8]
  PIN out0[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 496.890 516.985 497.170 520.985 ;
    END
  END out0[9]
  PIN out1[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 335.890 516.985 336.170 520.985 ;
    END
  END out1[0]
  PIN out1[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 355.000 510.265 355.600 ;
    END
  END out1[10]
  PIN out1[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 447.480 510.265 448.080 ;
    END
  END out1[11]
  PIN out1[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END out1[12]
  PIN out1[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END out1[13]
  PIN out1[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.170 516.985 45.450 520.985 ;
    END
  END out1[14]
  PIN out1[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 315.650 516.985 315.930 520.985 ;
    END
  END out1[15]
  PIN out1[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END out1[16]
  PIN out1[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 193.160 510.265 193.760 ;
    END
  END out1[17]
  PIN out1[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.650 516.985 39.930 520.985 ;
    END
  END out1[18]
  PIN out1[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END out1[19]
  PIN out1[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END out1[1]
  PIN out1[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 485.560 510.265 486.160 ;
    END
  END out1[20]
  PIN out1[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 434.330 516.985 434.610 520.985 ;
    END
  END out1[21]
  PIN out1[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END out1[22]
  PIN out1[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END out1[23]
  PIN out1[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.490 516.985 133.770 520.985 ;
    END
  END out1[24]
  PIN out1[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END out1[25]
  PIN out1[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END out1[26]
  PIN out1[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 492.290 516.985 492.570 520.985 ;
    END
  END out1[27]
  PIN out1[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 170.040 510.265 170.640 ;
    END
  END out1[28]
  PIN out1[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END out1[29]
  PIN out1[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END out1[2]
  PIN out1[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END out1[30]
  PIN out1[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 516.985 14.170 520.985 ;
    END
  END out1[31]
  PIN out1[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 70.760 510.265 71.360 ;
    END
  END out1[3]
  PIN out1[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END out1[4]
  PIN out1[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END out1[5]
  PIN out1[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END out1[6]
  PIN out1[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 186.360 510.265 186.960 ;
    END
  END out1[7]
  PIN out1[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 221.810 516.985 222.090 520.985 ;
    END
  END out1[8]
  PIN out1[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.010 516.985 139.290 520.985 ;
    END
  END out1[9]
  PIN out2[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END out2[0]
  PIN out2[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END out2[10]
  PIN out2[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 516.985 102.490 520.985 ;
    END
  END out2[11]
  PIN out2[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 140.120 510.265 140.720 ;
    END
  END out2[12]
  PIN out2[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END out2[13]
  PIN out2[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END out2[14]
  PIN out2[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 253.090 516.985 253.370 520.985 ;
    END
  END out2[15]
  PIN out2[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 320.250 516.985 320.530 520.985 ;
    END
  END out2[16]
  PIN out2[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 4.000 ;
    END
  END out2[17]
  PIN out2[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 401.240 510.265 401.840 ;
    END
  END out2[18]
  PIN out2[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END out2[19]
  PIN out2[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END out2[1]
  PIN out2[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 154.650 516.985 154.930 520.985 ;
    END
  END out2[20]
  PIN out2[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END out2[21]
  PIN out2[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 508.680 510.265 509.280 ;
    END
  END out2[22]
  PIN out2[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END out2[23]
  PIN out2[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 239.400 510.265 240.000 ;
    END
  END out2[24]
  PIN out2[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END out2[25]
  PIN out2[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 47.640 510.265 48.240 ;
    END
  END out2[26]
  PIN out2[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END out2[27]
  PIN out2[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 455.490 516.985 455.770 520.985 ;
    END
  END out2[28]
  PIN out2[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END out2[29]
  PIN out2[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 247.570 516.985 247.850 520.985 ;
    END
  END out2[2]
  PIN out2[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END out2[30]
  PIN out2[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END out2[31]
  PIN out2[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.330 516.985 66.610 520.985 ;
    END
  END out2[3]
  PIN out2[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 403.970 516.985 404.250 520.985 ;
    END
  END out2[4]
  PIN out2[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.050 516.985 196.330 520.985 ;
    END
  END out2[5]
  PIN out2[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END out2[6]
  PIN out2[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 200.650 516.985 200.930 520.985 ;
    END
  END out2[7]
  PIN out2[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END out2[8]
  PIN out2[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 62.600 510.265 63.200 ;
    END
  END out2[9]
  PIN out3[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END out3[0]
  PIN out3[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 449.970 516.985 450.250 520.985 ;
    END
  END out3[10]
  PIN out3[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 288.970 516.985 289.250 520.985 ;
    END
  END out3[11]
  PIN out3[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 361.650 516.985 361.930 520.985 ;
    END
  END out3[12]
  PIN out3[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END out3[13]
  PIN out3[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END out3[14]
  PIN out3[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 293.800 510.265 294.400 ;
    END
  END out3[15]
  PIN out3[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END out3[16]
  PIN out3[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END out3[17]
  PIN out3[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 372.690 516.985 372.970 520.985 ;
    END
  END out3[18]
  PIN out3[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 516.985 96.970 520.985 ;
    END
  END out3[19]
  PIN out3[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 516.985 61.090 520.985 ;
    END
  END out3[1]
  PIN out3[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END out3[20]
  PIN out3[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END out3[21]
  PIN out3[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END out3[22]
  PIN out3[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 273.330 516.985 273.610 520.985 ;
    END
  END out3[23]
  PIN out3[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END out3[24]
  PIN out3[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 85.720 510.265 86.320 ;
    END
  END out3[25]
  PIN out3[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END out3[26]
  PIN out3[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 516.985 8.650 520.985 ;
    END
  END out3[27]
  PIN out3[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 377.290 516.985 377.570 520.985 ;
    END
  END out3[28]
  PIN out3[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 419.610 516.985 419.890 520.985 ;
    END
  END out3[29]
  PIN out3[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END out3[2]
  PIN out3[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END out3[30]
  PIN out3[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END out3[31]
  PIN out3[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END out3[3]
  PIN out3[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END out3[4]
  PIN out3[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 237.450 516.985 237.730 520.985 ;
    END
  END out3[5]
  PIN out3[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END out3[6]
  PIN out3[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 506.265 9.560 510.265 10.160 ;
    END
  END out3[7]
  PIN out3[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END out3[8]
  PIN out3[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.410 516.985 502.690 520.985 ;
    END
  END out3[9]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END rst
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 504.620 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 504.620 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 504.620 508.725 ;
      LAYER met1 ;
        RECT 2.830 4.460 507.310 516.760 ;
      LAYER met2 ;
        RECT 2.860 516.705 3.490 516.985 ;
        RECT 4.330 516.705 8.090 516.985 ;
        RECT 8.930 516.705 13.610 516.985 ;
        RECT 14.450 516.705 19.130 516.985 ;
        RECT 19.970 516.705 23.730 516.985 ;
        RECT 24.570 516.705 29.250 516.985 ;
        RECT 30.090 516.705 34.770 516.985 ;
        RECT 35.610 516.705 39.370 516.985 ;
        RECT 40.210 516.705 44.890 516.985 ;
        RECT 45.730 516.705 50.410 516.985 ;
        RECT 51.250 516.705 55.010 516.985 ;
        RECT 55.850 516.705 60.530 516.985 ;
        RECT 61.370 516.705 66.050 516.985 ;
        RECT 66.890 516.705 70.650 516.985 ;
        RECT 71.490 516.705 76.170 516.985 ;
        RECT 77.010 516.705 80.770 516.985 ;
        RECT 81.610 516.705 86.290 516.985 ;
        RECT 87.130 516.705 91.810 516.985 ;
        RECT 92.650 516.705 96.410 516.985 ;
        RECT 97.250 516.705 101.930 516.985 ;
        RECT 102.770 516.705 107.450 516.985 ;
        RECT 108.290 516.705 112.050 516.985 ;
        RECT 112.890 516.705 117.570 516.985 ;
        RECT 118.410 516.705 123.090 516.985 ;
        RECT 123.930 516.705 127.690 516.985 ;
        RECT 128.530 516.705 133.210 516.985 ;
        RECT 134.050 516.705 138.730 516.985 ;
        RECT 139.570 516.705 143.330 516.985 ;
        RECT 144.170 516.705 148.850 516.985 ;
        RECT 149.690 516.705 154.370 516.985 ;
        RECT 155.210 516.705 158.970 516.985 ;
        RECT 159.810 516.705 164.490 516.985 ;
        RECT 165.330 516.705 169.090 516.985 ;
        RECT 169.930 516.705 174.610 516.985 ;
        RECT 175.450 516.705 180.130 516.985 ;
        RECT 180.970 516.705 184.730 516.985 ;
        RECT 185.570 516.705 190.250 516.985 ;
        RECT 191.090 516.705 195.770 516.985 ;
        RECT 196.610 516.705 200.370 516.985 ;
        RECT 201.210 516.705 205.890 516.985 ;
        RECT 206.730 516.705 211.410 516.985 ;
        RECT 212.250 516.705 216.010 516.985 ;
        RECT 216.850 516.705 221.530 516.985 ;
        RECT 222.370 516.705 227.050 516.985 ;
        RECT 227.890 516.705 231.650 516.985 ;
        RECT 232.490 516.705 237.170 516.985 ;
        RECT 238.010 516.705 242.690 516.985 ;
        RECT 243.530 516.705 247.290 516.985 ;
        RECT 248.130 516.705 252.810 516.985 ;
        RECT 253.650 516.705 257.410 516.985 ;
        RECT 258.250 516.705 262.930 516.985 ;
        RECT 263.770 516.705 268.450 516.985 ;
        RECT 269.290 516.705 273.050 516.985 ;
        RECT 273.890 516.705 278.570 516.985 ;
        RECT 279.410 516.705 284.090 516.985 ;
        RECT 284.930 516.705 288.690 516.985 ;
        RECT 289.530 516.705 294.210 516.985 ;
        RECT 295.050 516.705 299.730 516.985 ;
        RECT 300.570 516.705 304.330 516.985 ;
        RECT 305.170 516.705 309.850 516.985 ;
        RECT 310.690 516.705 315.370 516.985 ;
        RECT 316.210 516.705 319.970 516.985 ;
        RECT 320.810 516.705 325.490 516.985 ;
        RECT 326.330 516.705 331.010 516.985 ;
        RECT 331.850 516.705 335.610 516.985 ;
        RECT 336.450 516.705 341.130 516.985 ;
        RECT 341.970 516.705 345.730 516.985 ;
        RECT 346.570 516.705 351.250 516.985 ;
        RECT 352.090 516.705 356.770 516.985 ;
        RECT 357.610 516.705 361.370 516.985 ;
        RECT 362.210 516.705 366.890 516.985 ;
        RECT 367.730 516.705 372.410 516.985 ;
        RECT 373.250 516.705 377.010 516.985 ;
        RECT 377.850 516.705 382.530 516.985 ;
        RECT 383.370 516.705 388.050 516.985 ;
        RECT 388.890 516.705 392.650 516.985 ;
        RECT 393.490 516.705 398.170 516.985 ;
        RECT 399.010 516.705 403.690 516.985 ;
        RECT 404.530 516.705 408.290 516.985 ;
        RECT 409.130 516.705 413.810 516.985 ;
        RECT 414.650 516.705 419.330 516.985 ;
        RECT 420.170 516.705 423.930 516.985 ;
        RECT 424.770 516.705 429.450 516.985 ;
        RECT 430.290 516.705 434.050 516.985 ;
        RECT 434.890 516.705 439.570 516.985 ;
        RECT 440.410 516.705 445.090 516.985 ;
        RECT 445.930 516.705 449.690 516.985 ;
        RECT 450.530 516.705 455.210 516.985 ;
        RECT 456.050 516.705 460.730 516.985 ;
        RECT 461.570 516.705 465.330 516.985 ;
        RECT 466.170 516.705 470.850 516.985 ;
        RECT 471.690 516.705 476.370 516.985 ;
        RECT 477.210 516.705 480.970 516.985 ;
        RECT 481.810 516.705 486.490 516.985 ;
        RECT 487.330 516.705 492.010 516.985 ;
        RECT 492.850 516.705 496.610 516.985 ;
        RECT 497.450 516.705 502.130 516.985 ;
        RECT 502.970 516.705 506.730 516.985 ;
        RECT 2.860 4.280 507.280 516.705 ;
        RECT 3.410 4.000 7.170 4.280 ;
        RECT 8.010 4.000 12.690 4.280 ;
        RECT 13.530 4.000 17.290 4.280 ;
        RECT 18.130 4.000 22.810 4.280 ;
        RECT 23.650 4.000 28.330 4.280 ;
        RECT 29.170 4.000 32.930 4.280 ;
        RECT 33.770 4.000 38.450 4.280 ;
        RECT 39.290 4.000 43.970 4.280 ;
        RECT 44.810 4.000 48.570 4.280 ;
        RECT 49.410 4.000 54.090 4.280 ;
        RECT 54.930 4.000 59.610 4.280 ;
        RECT 60.450 4.000 64.210 4.280 ;
        RECT 65.050 4.000 69.730 4.280 ;
        RECT 70.570 4.000 75.250 4.280 ;
        RECT 76.090 4.000 79.850 4.280 ;
        RECT 80.690 4.000 85.370 4.280 ;
        RECT 86.210 4.000 89.970 4.280 ;
        RECT 90.810 4.000 95.490 4.280 ;
        RECT 96.330 4.000 101.010 4.280 ;
        RECT 101.850 4.000 105.610 4.280 ;
        RECT 106.450 4.000 111.130 4.280 ;
        RECT 111.970 4.000 116.650 4.280 ;
        RECT 117.490 4.000 121.250 4.280 ;
        RECT 122.090 4.000 126.770 4.280 ;
        RECT 127.610 4.000 132.290 4.280 ;
        RECT 133.130 4.000 136.890 4.280 ;
        RECT 137.730 4.000 142.410 4.280 ;
        RECT 143.250 4.000 147.930 4.280 ;
        RECT 148.770 4.000 152.530 4.280 ;
        RECT 153.370 4.000 158.050 4.280 ;
        RECT 158.890 4.000 163.570 4.280 ;
        RECT 164.410 4.000 168.170 4.280 ;
        RECT 169.010 4.000 173.690 4.280 ;
        RECT 174.530 4.000 178.290 4.280 ;
        RECT 179.130 4.000 183.810 4.280 ;
        RECT 184.650 4.000 189.330 4.280 ;
        RECT 190.170 4.000 193.930 4.280 ;
        RECT 194.770 4.000 199.450 4.280 ;
        RECT 200.290 4.000 204.970 4.280 ;
        RECT 205.810 4.000 209.570 4.280 ;
        RECT 210.410 4.000 215.090 4.280 ;
        RECT 215.930 4.000 220.610 4.280 ;
        RECT 221.450 4.000 225.210 4.280 ;
        RECT 226.050 4.000 230.730 4.280 ;
        RECT 231.570 4.000 236.250 4.280 ;
        RECT 237.090 4.000 240.850 4.280 ;
        RECT 241.690 4.000 246.370 4.280 ;
        RECT 247.210 4.000 251.890 4.280 ;
        RECT 252.730 4.000 256.490 4.280 ;
        RECT 257.330 4.000 262.010 4.280 ;
        RECT 262.850 4.000 266.610 4.280 ;
        RECT 267.450 4.000 272.130 4.280 ;
        RECT 272.970 4.000 277.650 4.280 ;
        RECT 278.490 4.000 282.250 4.280 ;
        RECT 283.090 4.000 287.770 4.280 ;
        RECT 288.610 4.000 293.290 4.280 ;
        RECT 294.130 4.000 297.890 4.280 ;
        RECT 298.730 4.000 303.410 4.280 ;
        RECT 304.250 4.000 308.930 4.280 ;
        RECT 309.770 4.000 313.530 4.280 ;
        RECT 314.370 4.000 319.050 4.280 ;
        RECT 319.890 4.000 324.570 4.280 ;
        RECT 325.410 4.000 329.170 4.280 ;
        RECT 330.010 4.000 334.690 4.280 ;
        RECT 335.530 4.000 340.210 4.280 ;
        RECT 341.050 4.000 344.810 4.280 ;
        RECT 345.650 4.000 350.330 4.280 ;
        RECT 351.170 4.000 354.930 4.280 ;
        RECT 355.770 4.000 360.450 4.280 ;
        RECT 361.290 4.000 365.970 4.280 ;
        RECT 366.810 4.000 370.570 4.280 ;
        RECT 371.410 4.000 376.090 4.280 ;
        RECT 376.930 4.000 381.610 4.280 ;
        RECT 382.450 4.000 386.210 4.280 ;
        RECT 387.050 4.000 391.730 4.280 ;
        RECT 392.570 4.000 397.250 4.280 ;
        RECT 398.090 4.000 401.850 4.280 ;
        RECT 402.690 4.000 407.370 4.280 ;
        RECT 408.210 4.000 412.890 4.280 ;
        RECT 413.730 4.000 417.490 4.280 ;
        RECT 418.330 4.000 423.010 4.280 ;
        RECT 423.850 4.000 428.530 4.280 ;
        RECT 429.370 4.000 433.130 4.280 ;
        RECT 433.970 4.000 438.650 4.280 ;
        RECT 439.490 4.000 443.250 4.280 ;
        RECT 444.090 4.000 448.770 4.280 ;
        RECT 449.610 4.000 454.290 4.280 ;
        RECT 455.130 4.000 458.890 4.280 ;
        RECT 459.730 4.000 464.410 4.280 ;
        RECT 465.250 4.000 469.930 4.280 ;
        RECT 470.770 4.000 474.530 4.280 ;
        RECT 475.370 4.000 480.050 4.280 ;
        RECT 480.890 4.000 485.570 4.280 ;
        RECT 486.410 4.000 490.170 4.280 ;
        RECT 491.010 4.000 495.690 4.280 ;
        RECT 496.530 4.000 501.210 4.280 ;
        RECT 502.050 4.000 505.810 4.280 ;
        RECT 506.650 4.000 507.280 4.280 ;
      LAYER met3 ;
        RECT 4.400 509.680 506.265 510.505 ;
        RECT 4.400 509.640 505.865 509.680 ;
        RECT 4.000 508.280 505.865 509.640 ;
        RECT 4.000 504.240 506.265 508.280 ;
        RECT 4.400 502.840 506.265 504.240 ;
        RECT 4.000 501.520 506.265 502.840 ;
        RECT 4.000 500.120 505.865 501.520 ;
        RECT 4.000 496.080 506.265 500.120 ;
        RECT 4.400 494.720 506.265 496.080 ;
        RECT 4.400 494.680 505.865 494.720 ;
        RECT 4.000 493.320 505.865 494.680 ;
        RECT 4.000 487.920 506.265 493.320 ;
        RECT 4.400 486.560 506.265 487.920 ;
        RECT 4.400 486.520 505.865 486.560 ;
        RECT 4.000 485.160 505.865 486.520 ;
        RECT 4.000 481.120 506.265 485.160 ;
        RECT 4.400 479.720 506.265 481.120 ;
        RECT 4.000 478.400 506.265 479.720 ;
        RECT 4.000 477.000 505.865 478.400 ;
        RECT 4.000 472.960 506.265 477.000 ;
        RECT 4.400 471.600 506.265 472.960 ;
        RECT 4.400 471.560 505.865 471.600 ;
        RECT 4.000 470.200 505.865 471.560 ;
        RECT 4.000 464.800 506.265 470.200 ;
        RECT 4.400 463.440 506.265 464.800 ;
        RECT 4.400 463.400 505.865 463.440 ;
        RECT 4.000 462.040 505.865 463.400 ;
        RECT 4.000 458.000 506.265 462.040 ;
        RECT 4.400 456.600 506.265 458.000 ;
        RECT 4.000 455.280 506.265 456.600 ;
        RECT 4.000 453.880 505.865 455.280 ;
        RECT 4.000 449.840 506.265 453.880 ;
        RECT 4.400 448.480 506.265 449.840 ;
        RECT 4.400 448.440 505.865 448.480 ;
        RECT 4.000 447.080 505.865 448.440 ;
        RECT 4.000 441.680 506.265 447.080 ;
        RECT 4.400 440.320 506.265 441.680 ;
        RECT 4.400 440.280 505.865 440.320 ;
        RECT 4.000 438.920 505.865 440.280 ;
        RECT 4.000 434.880 506.265 438.920 ;
        RECT 4.400 433.480 506.265 434.880 ;
        RECT 4.000 432.160 506.265 433.480 ;
        RECT 4.000 430.760 505.865 432.160 ;
        RECT 4.000 426.720 506.265 430.760 ;
        RECT 4.400 425.360 506.265 426.720 ;
        RECT 4.400 425.320 505.865 425.360 ;
        RECT 4.000 423.960 505.865 425.320 ;
        RECT 4.000 418.560 506.265 423.960 ;
        RECT 4.400 417.200 506.265 418.560 ;
        RECT 4.400 417.160 505.865 417.200 ;
        RECT 4.000 415.800 505.865 417.160 ;
        RECT 4.000 411.760 506.265 415.800 ;
        RECT 4.400 410.360 506.265 411.760 ;
        RECT 4.000 409.040 506.265 410.360 ;
        RECT 4.000 407.640 505.865 409.040 ;
        RECT 4.000 403.600 506.265 407.640 ;
        RECT 4.400 402.240 506.265 403.600 ;
        RECT 4.400 402.200 505.865 402.240 ;
        RECT 4.000 400.840 505.865 402.200 ;
        RECT 4.000 395.440 506.265 400.840 ;
        RECT 4.400 394.080 506.265 395.440 ;
        RECT 4.400 394.040 505.865 394.080 ;
        RECT 4.000 392.680 505.865 394.040 ;
        RECT 4.000 388.640 506.265 392.680 ;
        RECT 4.400 387.280 506.265 388.640 ;
        RECT 4.400 387.240 505.865 387.280 ;
        RECT 4.000 385.880 505.865 387.240 ;
        RECT 4.000 380.480 506.265 385.880 ;
        RECT 4.400 379.120 506.265 380.480 ;
        RECT 4.400 379.080 505.865 379.120 ;
        RECT 4.000 377.720 505.865 379.080 ;
        RECT 4.000 373.680 506.265 377.720 ;
        RECT 4.400 372.280 506.265 373.680 ;
        RECT 4.000 370.960 506.265 372.280 ;
        RECT 4.000 369.560 505.865 370.960 ;
        RECT 4.000 365.520 506.265 369.560 ;
        RECT 4.400 364.160 506.265 365.520 ;
        RECT 4.400 364.120 505.865 364.160 ;
        RECT 4.000 362.760 505.865 364.120 ;
        RECT 4.000 357.360 506.265 362.760 ;
        RECT 4.400 356.000 506.265 357.360 ;
        RECT 4.400 355.960 505.865 356.000 ;
        RECT 4.000 354.600 505.865 355.960 ;
        RECT 4.000 350.560 506.265 354.600 ;
        RECT 4.400 349.160 506.265 350.560 ;
        RECT 4.000 347.840 506.265 349.160 ;
        RECT 4.000 346.440 505.865 347.840 ;
        RECT 4.000 342.400 506.265 346.440 ;
        RECT 4.400 341.040 506.265 342.400 ;
        RECT 4.400 341.000 505.865 341.040 ;
        RECT 4.000 339.640 505.865 341.000 ;
        RECT 4.000 334.240 506.265 339.640 ;
        RECT 4.400 332.880 506.265 334.240 ;
        RECT 4.400 332.840 505.865 332.880 ;
        RECT 4.000 331.480 505.865 332.840 ;
        RECT 4.000 327.440 506.265 331.480 ;
        RECT 4.400 326.040 506.265 327.440 ;
        RECT 4.000 324.720 506.265 326.040 ;
        RECT 4.000 323.320 505.865 324.720 ;
        RECT 4.000 319.280 506.265 323.320 ;
        RECT 4.400 317.920 506.265 319.280 ;
        RECT 4.400 317.880 505.865 317.920 ;
        RECT 4.000 316.520 505.865 317.880 ;
        RECT 4.000 311.120 506.265 316.520 ;
        RECT 4.400 309.760 506.265 311.120 ;
        RECT 4.400 309.720 505.865 309.760 ;
        RECT 4.000 308.360 505.865 309.720 ;
        RECT 4.000 304.320 506.265 308.360 ;
        RECT 4.400 302.920 506.265 304.320 ;
        RECT 4.000 301.600 506.265 302.920 ;
        RECT 4.000 300.200 505.865 301.600 ;
        RECT 4.000 296.160 506.265 300.200 ;
        RECT 4.400 294.800 506.265 296.160 ;
        RECT 4.400 294.760 505.865 294.800 ;
        RECT 4.000 293.400 505.865 294.760 ;
        RECT 4.000 288.000 506.265 293.400 ;
        RECT 4.400 286.640 506.265 288.000 ;
        RECT 4.400 286.600 505.865 286.640 ;
        RECT 4.000 285.240 505.865 286.600 ;
        RECT 4.000 281.200 506.265 285.240 ;
        RECT 4.400 279.800 506.265 281.200 ;
        RECT 4.000 278.480 506.265 279.800 ;
        RECT 4.000 277.080 505.865 278.480 ;
        RECT 4.000 273.040 506.265 277.080 ;
        RECT 4.400 271.680 506.265 273.040 ;
        RECT 4.400 271.640 505.865 271.680 ;
        RECT 4.000 270.280 505.865 271.640 ;
        RECT 4.000 264.880 506.265 270.280 ;
        RECT 4.400 263.520 506.265 264.880 ;
        RECT 4.400 263.480 505.865 263.520 ;
        RECT 4.000 262.120 505.865 263.480 ;
        RECT 4.000 258.080 506.265 262.120 ;
        RECT 4.400 256.720 506.265 258.080 ;
        RECT 4.400 256.680 505.865 256.720 ;
        RECT 4.000 255.320 505.865 256.680 ;
        RECT 4.000 249.920 506.265 255.320 ;
        RECT 4.400 248.560 506.265 249.920 ;
        RECT 4.400 248.520 505.865 248.560 ;
        RECT 4.000 247.160 505.865 248.520 ;
        RECT 4.000 243.120 506.265 247.160 ;
        RECT 4.400 241.720 506.265 243.120 ;
        RECT 4.000 240.400 506.265 241.720 ;
        RECT 4.000 239.000 505.865 240.400 ;
        RECT 4.000 234.960 506.265 239.000 ;
        RECT 4.400 233.600 506.265 234.960 ;
        RECT 4.400 233.560 505.865 233.600 ;
        RECT 4.000 232.200 505.865 233.560 ;
        RECT 4.000 226.800 506.265 232.200 ;
        RECT 4.400 225.440 506.265 226.800 ;
        RECT 4.400 225.400 505.865 225.440 ;
        RECT 4.000 224.040 505.865 225.400 ;
        RECT 4.000 220.000 506.265 224.040 ;
        RECT 4.400 218.600 506.265 220.000 ;
        RECT 4.000 217.280 506.265 218.600 ;
        RECT 4.000 215.880 505.865 217.280 ;
        RECT 4.000 211.840 506.265 215.880 ;
        RECT 4.400 210.480 506.265 211.840 ;
        RECT 4.400 210.440 505.865 210.480 ;
        RECT 4.000 209.080 505.865 210.440 ;
        RECT 4.000 203.680 506.265 209.080 ;
        RECT 4.400 202.320 506.265 203.680 ;
        RECT 4.400 202.280 505.865 202.320 ;
        RECT 4.000 200.920 505.865 202.280 ;
        RECT 4.000 196.880 506.265 200.920 ;
        RECT 4.400 195.480 506.265 196.880 ;
        RECT 4.000 194.160 506.265 195.480 ;
        RECT 4.000 192.760 505.865 194.160 ;
        RECT 4.000 188.720 506.265 192.760 ;
        RECT 4.400 187.360 506.265 188.720 ;
        RECT 4.400 187.320 505.865 187.360 ;
        RECT 4.000 185.960 505.865 187.320 ;
        RECT 4.000 180.560 506.265 185.960 ;
        RECT 4.400 179.200 506.265 180.560 ;
        RECT 4.400 179.160 505.865 179.200 ;
        RECT 4.000 177.800 505.865 179.160 ;
        RECT 4.000 173.760 506.265 177.800 ;
        RECT 4.400 172.360 506.265 173.760 ;
        RECT 4.000 171.040 506.265 172.360 ;
        RECT 4.000 169.640 505.865 171.040 ;
        RECT 4.000 165.600 506.265 169.640 ;
        RECT 4.400 164.240 506.265 165.600 ;
        RECT 4.400 164.200 505.865 164.240 ;
        RECT 4.000 162.840 505.865 164.200 ;
        RECT 4.000 157.440 506.265 162.840 ;
        RECT 4.400 156.080 506.265 157.440 ;
        RECT 4.400 156.040 505.865 156.080 ;
        RECT 4.000 154.680 505.865 156.040 ;
        RECT 4.000 150.640 506.265 154.680 ;
        RECT 4.400 149.240 506.265 150.640 ;
        RECT 4.000 147.920 506.265 149.240 ;
        RECT 4.000 146.520 505.865 147.920 ;
        RECT 4.000 142.480 506.265 146.520 ;
        RECT 4.400 141.120 506.265 142.480 ;
        RECT 4.400 141.080 505.865 141.120 ;
        RECT 4.000 139.720 505.865 141.080 ;
        RECT 4.000 134.320 506.265 139.720 ;
        RECT 4.400 132.960 506.265 134.320 ;
        RECT 4.400 132.920 505.865 132.960 ;
        RECT 4.000 131.560 505.865 132.920 ;
        RECT 4.000 127.520 506.265 131.560 ;
        RECT 4.400 126.160 506.265 127.520 ;
        RECT 4.400 126.120 505.865 126.160 ;
        RECT 4.000 124.760 505.865 126.120 ;
        RECT 4.000 119.360 506.265 124.760 ;
        RECT 4.400 118.000 506.265 119.360 ;
        RECT 4.400 117.960 505.865 118.000 ;
        RECT 4.000 116.600 505.865 117.960 ;
        RECT 4.000 112.560 506.265 116.600 ;
        RECT 4.400 111.160 506.265 112.560 ;
        RECT 4.000 109.840 506.265 111.160 ;
        RECT 4.000 108.440 505.865 109.840 ;
        RECT 4.000 104.400 506.265 108.440 ;
        RECT 4.400 103.040 506.265 104.400 ;
        RECT 4.400 103.000 505.865 103.040 ;
        RECT 4.000 101.640 505.865 103.000 ;
        RECT 4.000 96.240 506.265 101.640 ;
        RECT 4.400 94.880 506.265 96.240 ;
        RECT 4.400 94.840 505.865 94.880 ;
        RECT 4.000 93.480 505.865 94.840 ;
        RECT 4.000 89.440 506.265 93.480 ;
        RECT 4.400 88.040 506.265 89.440 ;
        RECT 4.000 86.720 506.265 88.040 ;
        RECT 4.000 85.320 505.865 86.720 ;
        RECT 4.000 81.280 506.265 85.320 ;
        RECT 4.400 79.920 506.265 81.280 ;
        RECT 4.400 79.880 505.865 79.920 ;
        RECT 4.000 78.520 505.865 79.880 ;
        RECT 4.000 73.120 506.265 78.520 ;
        RECT 4.400 71.760 506.265 73.120 ;
        RECT 4.400 71.720 505.865 71.760 ;
        RECT 4.000 70.360 505.865 71.720 ;
        RECT 4.000 66.320 506.265 70.360 ;
        RECT 4.400 64.920 506.265 66.320 ;
        RECT 4.000 63.600 506.265 64.920 ;
        RECT 4.000 62.200 505.865 63.600 ;
        RECT 4.000 58.160 506.265 62.200 ;
        RECT 4.400 56.800 506.265 58.160 ;
        RECT 4.400 56.760 505.865 56.800 ;
        RECT 4.000 55.400 505.865 56.760 ;
        RECT 4.000 50.000 506.265 55.400 ;
        RECT 4.400 48.640 506.265 50.000 ;
        RECT 4.400 48.600 505.865 48.640 ;
        RECT 4.000 47.240 505.865 48.600 ;
        RECT 4.000 43.200 506.265 47.240 ;
        RECT 4.400 41.800 506.265 43.200 ;
        RECT 4.000 40.480 506.265 41.800 ;
        RECT 4.000 39.080 505.865 40.480 ;
        RECT 4.000 35.040 506.265 39.080 ;
        RECT 4.400 33.680 506.265 35.040 ;
        RECT 4.400 33.640 505.865 33.680 ;
        RECT 4.000 32.280 505.865 33.640 ;
        RECT 4.000 26.880 506.265 32.280 ;
        RECT 4.400 25.520 506.265 26.880 ;
        RECT 4.400 25.480 505.865 25.520 ;
        RECT 4.000 24.120 505.865 25.480 ;
        RECT 4.000 20.080 506.265 24.120 ;
        RECT 4.400 18.680 506.265 20.080 ;
        RECT 4.000 17.360 506.265 18.680 ;
        RECT 4.000 15.960 505.865 17.360 ;
        RECT 4.000 11.920 506.265 15.960 ;
        RECT 4.400 10.560 506.265 11.920 ;
        RECT 4.400 10.520 505.865 10.560 ;
        RECT 4.000 9.160 505.865 10.520 ;
        RECT 4.000 4.255 506.265 9.160 ;
      LAYER met4 ;
        RECT 15.935 10.640 490.065 508.880 ;
      LAYER met5 ;
        RECT 5.520 179.670 504.620 487.630 ;
  END
END mac_cluster
END LIBRARY

